// Note: The license below is based on the template at:
// http://opensource.org/licenses/BSD-3-Clause
// Copyright (C) 2020 Regents of the University of Texas
//All rights reserved.

// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are
// met:

// o Redistributions of source code must retain the above copyright
//   notice, this list of conditions and the following disclaimer.

// o Redistributions in binary form must reproduce the above copyright
//   notice, this list of conditions and the following disclaimer in the
//   documentation and/or other materials provided with the distribution.

// o Neither the name of the copyright holders nor the names of its
//   contributors may be used to endorse or promote products derived
//   from this software without specific prior written permission.

// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
// A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT
// HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
// SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT
// LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
// DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
// THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

// Original Author(s):
// Mertcan Temel         <mert@utexas.edu>

// DO NOT REMOVE:
// This file is generated by Temel's multiplier generator. Download from https://github.com/temelmertcan/multgen.


// Specification module to help understand what the design implements.
module Merged_c42_SB4_JSkCond_16x16_14to0_spec (
        input logic [15:0] IN1,
        input logic [15:0] IN2,
        input logic [0:0] IN3, //redundant
        output logic design_is_correct, // is set to 1 iff the output of Merged_c42_SB4_JSkCond_16x16_14to0  matches its spec.
        output logic [14:0] design_res,
        output logic [14:0] spec_res);
    
    assign spec_res = signed'(IN1) * signed'(IN2) ;
    Merged_c42_SB4_JSkCond_16x16_14to0 mult(IN1, IN2, design_res);
    assign design_is_correct = ((spec_res == design_res) ? 1 : 0);
    
endmodule



module c42_SB4_9x9(
        input logic [8:0] IN1,
        input logic [8:0] IN2,
        output logic [14:0] result0,
        output logic [14:0] result1);
    
    
// Creating Partial Products 

    wire [8:0] mult = IN1;
    wire [8:0] mcand = IN2;
    wire [9:0] mcand_1x;
    wire [9:0] mcand_2x;
    assign mcand_1x = {{1{mcand[8]}},  mcand};
    assign mcand_2x = {{0{mcand[8]}},  mcand, 1'b0};
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[1] mult[0] 1'b0
    wire logic select_0_0, select_e_0, select_2x_0, tcomp0, select_ne_0, select_n2x_0;
    assign select_0_0 =  &{mult[1], mult[0], 1'b0} | ~|{mult[1], mult[0], 1'b0};
    assign select_e_0 = ((~ mult[1]) & (mult[0] ^ 1'b0));
    assign select_ne_0 = mult[1] &  (mult[0] ^ 1'b0);
    assign select_2x_0 = (~ mult[1]) & mult[0] & 1'b0;
    assign select_n2x_0 = mult[1] & (~ mult[0]) & (~ 1'b0);
    reg [9:0] pp_0;
    always @(*) begin
       case (1'b1)
          select_0_0   : pp_0 = 0; 
          select_e_0   : pp_0 = mcand_1x; 
          select_2x_0  : pp_0 = mcand_2x; 
          select_n2x_0 : pp_0 = (~ mcand_2x); 
          select_ne_0  : pp_0 = (~ mcand_1x); 
       endcase 
       pp_0[9] = ~pp_0[9]; // flip the MSB 
    end
    assign tcomp0 =  select_n2x_0 | select_ne_0;
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[3] mult[2] mult[1]
    wire logic select_0_1, select_e_1, select_2x_1, tcomp1, select_ne_1, select_n2x_1;
    assign select_0_1 =  &{mult[3], mult[2], mult[1]} | ~|{mult[3], mult[2], mult[1]};
    assign select_e_1 = ((~ mult[3]) & (mult[2] ^ mult[1]));
    assign select_ne_1 = mult[3] &  (mult[2] ^ mult[1]);
    assign select_2x_1 = (~ mult[3]) & mult[2] & mult[1];
    assign select_n2x_1 = mult[3] & (~ mult[2]) & (~ mult[1]);
    reg [9:0] pp_1;
    always @(*) begin
       case (1'b1)
          select_0_1   : pp_1 = 0; 
          select_e_1   : pp_1 = mcand_1x; 
          select_2x_1  : pp_1 = mcand_2x; 
          select_n2x_1 : pp_1 = (~ mcand_2x); 
          select_ne_1  : pp_1 = (~ mcand_1x); 
       endcase 
       pp_1[9] = ~pp_1[9]; // flip the MSB 
    end
    assign tcomp1 =  select_n2x_1 | select_ne_1;
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[5] mult[4] mult[3]
    wire logic select_0_2, select_e_2, select_2x_2, tcomp2, select_ne_2, select_n2x_2;
    assign select_0_2 =  &{mult[5], mult[4], mult[3]} | ~|{mult[5], mult[4], mult[3]};
    assign select_e_2 = ((~ mult[5]) & (mult[4] ^ mult[3]));
    assign select_ne_2 = mult[5] &  (mult[4] ^ mult[3]);
    assign select_2x_2 = (~ mult[5]) & mult[4] & mult[3];
    assign select_n2x_2 = mult[5] & (~ mult[4]) & (~ mult[3]);
    reg [9:0] pp_2;
    always @(*) begin
       case (1'b1)
          select_0_2   : pp_2 = 0; 
          select_e_2   : pp_2 = mcand_1x; 
          select_2x_2  : pp_2 = mcand_2x; 
          select_n2x_2 : pp_2 = (~ mcand_2x); 
          select_ne_2  : pp_2 = (~ mcand_1x); 
       endcase 
       pp_2[9] = ~pp_2[9]; // flip the MSB 
    end
    assign tcomp2 =  select_n2x_2 | select_ne_2;
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[7] mult[6] mult[5]
    wire logic select_0_3, select_e_3, select_2x_3, tcomp3, select_ne_3, select_n2x_3;
    assign select_0_3 =  &{mult[7], mult[6], mult[5]} | ~|{mult[7], mult[6], mult[5]};
    assign select_e_3 = ((~ mult[7]) & (mult[6] ^ mult[5]));
    assign select_ne_3 = mult[7] &  (mult[6] ^ mult[5]);
    assign select_2x_3 = (~ mult[7]) & mult[6] & mult[5];
    assign select_n2x_3 = mult[7] & (~ mult[6]) & (~ mult[5]);
    reg [9:0] pp_3;
    always @(*) begin
       case (1'b1)
          select_0_3   : pp_3 = 0; 
          select_e_3   : pp_3 = mcand_1x; 
          select_2x_3  : pp_3 = mcand_2x; 
          select_n2x_3 : pp_3 = (~ mcand_2x); 
          select_ne_3  : pp_3 = (~ mcand_1x); 
       endcase 
       pp_3[9] = ~pp_3[9]; // flip the MSB 
    end
    assign tcomp3 =  select_n2x_3 | select_ne_3;
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[8] mult[8] mult[7]
    wire logic select_0_4, select_e_4, select_2x_4, tcomp4, select_ne_4, select_n2x_4;
    assign select_0_4 =  &{mult[8], mult[8], mult[7]} | ~|{mult[8], mult[8], mult[7]};
    assign select_e_4 = ((~ mult[8]) & (mult[8] ^ mult[7]));
    assign select_ne_4 = mult[8] &  (mult[8] ^ mult[7]);
    assign select_2x_4 = (~ mult[8]) & mult[8] & mult[7];
    assign select_n2x_4 = mult[8] & (~ mult[8]) & (~ mult[7]);
    reg [9:0] pp_4;
    always @(*) begin
       case (1'b1)
          select_0_4   : pp_4 = 0; 
          select_e_4   : pp_4 = mcand_1x; 
          select_2x_4  : pp_4 = mcand_2x; 
          select_n2x_4 : pp_4 = (~ mcand_2x); 
          select_ne_4  : pp_4 = (~ mcand_1x); 
       endcase 
       pp_4[9] = ~pp_4[9]; // flip the MSB 
    end
    assign tcomp4 =  select_n2x_4 | select_ne_4;
    
    // The values to be summed in the summation tree, from LSB (left) to MSB:
     // pp_0[0] pp_0[1] pp_0[2] pp_0[3] pp_0[4] pp_0[5] pp_0[6] pp_0[7] pp_0[8] pp_0[9]   --      --      --      --      --      --      --      --    
     //   --      --    pp_1[0] pp_1[1] pp_1[2] pp_1[3] pp_1[4] pp_1[5] pp_1[6] pp_1[7] pp_1[8] pp_1[9]   --      --      --      --      --      --    
     //   --      --      --      --    pp_2[0] pp_2[1] pp_2[2] pp_2[3] pp_2[4] pp_2[5] pp_2[6] pp_2[7] pp_2[8] pp_2[9]   --      --      --      --    
     //   --      --      --      --      --      --    pp_3[0] pp_3[1] pp_3[2] pp_3[3] pp_3[4] pp_3[5] pp_3[6] pp_3[7] pp_3[8] pp_3[9]   --      --    
     //   --      --      --      --      --      --      --      --    pp_4[0] pp_4[1] pp_4[2] pp_4[3] pp_4[4] pp_4[5] pp_4[6] pp_4[7] pp_4[8] pp_4[9] 
     // tcomp0    --    tcomp1    --    tcomp2    --    tcomp3    --    tcomp4    --      --      --      --      --      --      --      --      --    
     //   --      --      --      --      --      --      --      --      --      --      --      --      --      --      --      --      --      --    
    
// Creating Summation Tree 

    
    // 4to2 compressor tree Stage 1
    
    wire cout0;
    wire [8:0] sum0;
    wire [8:0] carry0;
    Four2Two #(9) cmp42_0(
            .in1({pp_3[8], pp_2[9:8], pp_1[9:8], pp_0[9:6]}),
            .in2({pp_4[6], pp_3[7:6], pp_2[7:6], pp_1[7:4]}),
            .in3({1'b0, pp_4[5:4], pp_3[5:4], pp_2[5:2]}),
            .in4({3'b0, pp_4[3:2], pp_3[3:0]}),
            .cin(tcomp3),
            .sum(sum0),
            .carry(carry0),
            .cout(cout0));
    
    wire cout1;
    wire [1:0] sum1;
    wire [1:0] carry1;
    Four2Two #(2) cmp42_1(
            .in1({pp_4[1:0]}),
            .in2({1'b0, tcomp4}),
            .in3({2'b0}),
            .in4({2'b0}),
            .cin(1'b0),
            .sum(sum1),
            .carry(carry1),
            .cout(cout1));
    
    // 4to2 compressor tree Stage 2
    
    wire cout2;
    wire [12:0] sum2;
    wire [12:0] carry2;
    Four2Two #(13) cmp42_2(
            .in1({carry0[7:0], sum0[0], pp_0[5:2]}),
            .in2({sum0[8:1], 1'b0, pp_1[3:0]}),
            .in3({4'b0, carry1[1:0], sum1[0], 2'b0, pp_2[1:0], 1'b0, tcomp1}),
            .in4({4'b0, cout1, sum1[1], 4'b0, tcomp2, 2'b0}),
            .cin(1'b0),
            .sum(sum2),
            .carry(carry2),
            .cout(cout2));
    
    
    assign result0[14:0] = {carry2[11], carry2[10], carry2[9], carry2[8], carry2[7], carry2[6], carry2[5], carry2[4], carry2[3], carry2[2], carry2[1], carry2[0], sum2[0], pp_0[1], pp_0[0] };
    assign result1[14:0] = {sum2[12], sum2[11], sum2[10], sum2[9], sum2[8], sum2[7], sum2[6], sum2[5], sum2[4], sum2[3], sum2[2], sum2[1], 1'b0, 1'b0, tcomp0 };
endmodule



module Merged_c42_SB4_JSkCond_16x16_14to0(
        input logic [15:0] IN1,
        input logic [15:0] IN2,
        output logic [14:0] result);
    wire logic [14:0] m1_0;
    wire logic [14:0] m1_1;
    wire logic [14:0] m2_0;
    wire logic [14:0] m2_1;
    wire logic [14:0] m3_0;
    wire logic [14:0] m3_1;
    wire logic [14:0] m4_0;
    wire logic [14:0] m4_1;
    
    c42_SB4_9x9 m1 ({1'b0, IN1[7:0]}, {1'b0, IN2[7:0]}, m1_0, m1_1);
    c42_SB4_9x9 m2 ({IN2[15], IN2[15:8]}, {1'b0, IN1[7:0]}, m2_0, m2_1);
    c42_SB4_9x9 m3 ({IN1[15], IN1[15:8]}, {1'b0, IN2[7:0]}, m3_0, m3_1);
    c42_SB4_9x9 m4 ({IN1[15],IN1[15:8]}, {IN2[15], IN2[15:8]}, m4_0, m4_1);
    
    
    // The values to be summed in the summation tree, from LSB (left) to MSB:
     // m1_0[0]  m1_0[1]  m1_0[2]  m1_0[3]  m1_0[4]  m1_0[5]  m1_0[6]  m1_0[7]  m1_0[8]  m1_0[9]  m1_0[10] m1_0[11] m1_0[12] m1_0[13] m1_0[14] 
     // m1_1[0]    --       --     m1_1[3]  m1_1[4]  m1_1[5]  m1_1[6]  m1_1[7]  m1_1[8]  m1_1[9]  m1_1[10] m1_1[11] m1_1[12] m1_1[13] m1_1[14] 
     //   --       --       --       --       --       --       --       --     m2_0[0]  m2_0[1]  m2_0[2]  m2_0[3]  m2_0[4]  m2_0[5]  m2_0[6]  
     //   --       --       --       --       --       --       --       --     m2_1[0]    --       --     m2_1[3]  m2_1[4]  m2_1[5]  m2_1[6]  
     //   --       --       --       --       --       --       --       --     m3_0[0]  m3_0[1]  m3_0[2]  m3_0[3]  m3_0[4]  m3_0[5]  m3_0[6]  
     //   --       --       --       --       --       --       --       --     m3_1[0]    --       --     m3_1[3]  m3_1[4]  m3_1[5]  m3_1[6]  
     //   --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --       --     1'b1     1'b1       --     1'b1       --     1'b1     
    
    // 4to2 compressor tree Stage 1
    
    wire cout0;
    wire [6:0] sum0;
    wire [6:0] carry0;
    Four2Two #(7) cmp42_0(
            .in1({m1_0[14:8]}),
            .in2({m1_1[14:8]}),
            .in3({m2_0[6:0]}),
            .in4({m2_1[6:3], m3_0[2:1], m2_1[0]}),
            .cin(m3_0[0]),
            .sum(sum0),
            .carry(carry0),
            .cout(cout0));
    
    wire cout1;
    wire [3:0] sum1;
    wire [3:0] carry1;
    Four2Two #(4) cmp42_1(
            .in1({m3_0[6:3]}),
            .in2({m3_1[6:3]}),
            .in3({1'b1, 1'b0, 1'b1, 1'b0}),
            .in4({4'b0}),
            .cin(1'b0),
            .sum(sum1),
            .carry(carry1),
            .cout(cout1));
    
    // 4to2 compressor tree Stage 2
    
    wire cout2;
    wire [5:0] sum2;
    wire [5:0] carry2;
    Four2Two #(6) cmp42_2(
            .in1({carry0[5:2], 1'b1, 1'b1}),
            .in2({sum0[6:3], carry0[1:0]}),
            .in3({carry1[2:0], sum1[0], sum0[2:1]}),
            .in4({sum1[3:1], 3'b0}),
            .cin(1'b0),
            .sum(sum2),
            .carry(carry2),
            .cout(cout2));
    
    logic [15:0] adder_result;
    JSkCond_15 final_adder ({carry2[4], carry2[3], carry2[2], carry2[1], carry2[0], sum2[0], m3_1[0], m1_0[7], m1_0[6], m1_0[5], m1_0[4], m1_0[3], m1_0[2], m1_0[1], m1_0[0] }, {sum2[5], sum2[4], sum2[3], sum2[2], sum2[1], 1'b0, sum0[0], m1_1[7], m1_1[6], m1_1[5], m1_1[4], m1_1[3], 1'b0, 1'b0, m1_1[0] }, adder_result );
    assign result[14:0] = adder_result[14:0];

endmodule

module JSkCond_15 ( 
        input logic [14:0] IN1,
        input logic [14:0] IN2,
        output logic [15:0] OUT);
    
    wire logic [14:0] p_0;
    wire logic [14:0] g_0;
    assign g_0 = IN1 & IN2;
    assign p_0 = IN1 ^ IN2;
    
    // J. Sklansky – Conditional Adder 

    
    // Stage 1 - prop from 1 to 1 per group.
    wire logic p_1_1;
    wire logic g_1_1;
    assign p_1_1 = p_0[1] & p_0[0];
    assign g_1_1 = (p_0[1] & g_0[0]) | g_0[1];
    wire logic p_1_3;
    wire logic g_1_3;
    assign p_1_3 = p_0[3] & p_0[2];
    assign g_1_3 = (p_0[3] & g_0[2]) | g_0[3];
    wire logic p_1_5;
    wire logic g_1_5;
    assign p_1_5 = p_0[5] & p_0[4];
    assign g_1_5 = (p_0[5] & g_0[4]) | g_0[5];
    wire logic p_1_7;
    wire logic g_1_7;
    assign p_1_7 = p_0[7] & p_0[6];
    assign g_1_7 = (p_0[7] & g_0[6]) | g_0[7];
    wire logic p_1_9;
    wire logic g_1_9;
    assign p_1_9 = p_0[9] & p_0[8];
    assign g_1_9 = (p_0[9] & g_0[8]) | g_0[9];
    wire logic p_1_11;
    wire logic g_1_11;
    assign p_1_11 = p_0[11] & p_0[10];
    assign g_1_11 = (p_0[11] & g_0[10]) | g_0[11];
    wire logic p_1_13;
    wire logic g_1_13;
    assign p_1_13 = p_0[13] & p_0[12];
    assign g_1_13 = (p_0[13] & g_0[12]) | g_0[13];
    
    // Stage 2 - prop from 1 to 2 per group.
    wire logic p_2_2;
    wire logic g_2_2;
    assign p_2_2 = p_0[2] & p_1_1;
    assign g_2_2 = (p_0[2] & g_1_1) | g_0[2];
    wire logic p_2_3;
    wire logic g_2_3;
    assign p_2_3 = p_1_3 & p_1_1;
    assign g_2_3 = (p_1_3 & g_1_1) | g_1_3;
    wire logic p_2_6;
    wire logic g_2_6;
    assign p_2_6 = p_0[6] & p_1_5;
    assign g_2_6 = (p_0[6] & g_1_5) | g_0[6];
    wire logic p_2_7;
    wire logic g_2_7;
    assign p_2_7 = p_1_7 & p_1_5;
    assign g_2_7 = (p_1_7 & g_1_5) | g_1_7;
    wire logic p_2_10;
    wire logic g_2_10;
    assign p_2_10 = p_0[10] & p_1_9;
    assign g_2_10 = (p_0[10] & g_1_9) | g_0[10];
    wire logic p_2_11;
    wire logic g_2_11;
    assign p_2_11 = p_1_11 & p_1_9;
    assign g_2_11 = (p_1_11 & g_1_9) | g_1_11;
    wire logic p_2_14;
    wire logic g_2_14;
    assign p_2_14 = p_0[14] & p_1_13;
    assign g_2_14 = (p_0[14] & g_1_13) | g_0[14];
    
    // Stage 3 - prop from 1 to 4 per group.
    wire logic p_3_4;
    wire logic g_3_4;
    assign p_3_4 = p_0[4] & p_2_3;
    assign g_3_4 = (p_0[4] & g_2_3) | g_0[4];
    wire logic p_3_5;
    wire logic g_3_5;
    assign p_3_5 = p_1_5 & p_2_3;
    assign g_3_5 = (p_1_5 & g_2_3) | g_1_5;
    wire logic p_3_6;
    wire logic g_3_6;
    assign p_3_6 = p_2_6 & p_2_3;
    assign g_3_6 = (p_2_6 & g_2_3) | g_2_6;
    wire logic p_3_7;
    wire logic g_3_7;
    assign p_3_7 = p_2_7 & p_2_3;
    assign g_3_7 = (p_2_7 & g_2_3) | g_2_7;
    wire logic p_3_12;
    wire logic g_3_12;
    assign p_3_12 = p_0[12] & p_2_11;
    assign g_3_12 = (p_0[12] & g_2_11) | g_0[12];
    wire logic p_3_13;
    wire logic g_3_13;
    assign p_3_13 = p_1_13 & p_2_11;
    assign g_3_13 = (p_1_13 & g_2_11) | g_1_13;
    wire logic p_3_14;
    wire logic g_3_14;
    assign p_3_14 = p_2_14 & p_2_11;
    assign g_3_14 = (p_2_14 & g_2_11) | g_2_14;
    
    // Stage 4 - prop from 1 to 8 per group.
    wire logic p_4_8;
    wire logic g_4_8;
    assign p_4_8 = p_0[8] & p_3_7;
    assign g_4_8 = (p_0[8] & g_3_7) | g_0[8];
    wire logic p_4_9;
    wire logic g_4_9;
    assign p_4_9 = p_1_9 & p_3_7;
    assign g_4_9 = (p_1_9 & g_3_7) | g_1_9;
    wire logic p_4_10;
    wire logic g_4_10;
    assign p_4_10 = p_2_10 & p_3_7;
    assign g_4_10 = (p_2_10 & g_3_7) | g_2_10;
    wire logic p_4_11;
    wire logic g_4_11;
    assign p_4_11 = p_2_11 & p_3_7;
    assign g_4_11 = (p_2_11 & g_3_7) | g_2_11;
    wire logic p_4_12;
    wire logic g_4_12;
    assign p_4_12 = p_3_12 & p_3_7;
    assign g_4_12 = (p_3_12 & g_3_7) | g_3_12;
    wire logic p_4_13;
    wire logic g_4_13;
    assign p_4_13 = p_3_13 & p_3_7;
    assign g_4_13 = (p_3_13 & g_3_7) | g_3_13;
    wire logic p_4_14;
    wire logic g_4_14;
    assign p_4_14 = p_3_14 & p_3_7;
    assign g_4_14 = (p_3_14 & g_3_7) | g_3_14;
    
    // JSkCondA postprocess 
    assign OUT[0] = p_0[0];
    assign OUT[1] = p_0[1] ^ g_0[0];
    assign OUT[2] = p_0[2] ^ g_1_1;
    assign OUT[3] = p_0[3] ^ g_2_2;
    assign OUT[4] = p_0[4] ^ g_2_3;
    assign OUT[5] = p_0[5] ^ g_3_4;
    assign OUT[6] = p_0[6] ^ g_3_5;
    assign OUT[7] = p_0[7] ^ g_3_6;
    assign OUT[8] = p_0[8] ^ g_3_7;
    assign OUT[9] = p_0[9] ^ g_4_8;
    assign OUT[10] = p_0[10] ^ g_4_9;
    assign OUT[11] = p_0[11] ^ g_4_10;
    assign OUT[12] = p_0[12] ^ g_4_11;
    assign OUT[13] = p_0[13] ^ g_4_12;
    assign OUT[14] = p_0[14] ^ g_4_13;
    assign OUT[15] = g_4_14;
endmodule

module JSkCond_15_spec (
        input logic [14:0] IN1,
        input logic [14:0] IN2,
        output logic adder_correct,
        output logic [15:0] spec_res);
    
    assign spec_res = IN1 + IN2;
    wire [15:0] adder_res;
    JSkCond_15 adder(IN1, IN2, adder_res);
    assign adder_correct = ((spec_res == adder_res) ? 1 : 0);
    
endmodule



module ha (
        input logic a,
        input logic b,
        output logic s,
        output logic c);
    
    assign s = a ^ b;
    assign c = a & b;
endmodule



module fa (
        input logic x,
        input logic y,
        input logic z,
        output logic s,
        output logic c);
    
    assign s = x ^ y ^ z;
    assign c = (x & y) | (x & z) | (y & z);
endmodule

module Four2Two 
        #(parameter WIDTH=1) (
        input logic [WIDTH-1:0] in1,
        input logic [WIDTH-1:0] in2,
        input logic [WIDTH-1:0] in3,
        input logic [WIDTH-1:0] in4,
        input logic cin,
        output logic [WIDTH-1:0] sum,
        output logic [WIDTH-1:0] carry,
        output logic cout);
    
    wire logic [WIDTH:0] temp1;
    assign temp1 = {((in1 ^ in2)&in3 | in1 & ~(in1^in2)),cin};
    assign sum = ((in1 ^ in2) ^ in3 ^ in4) ^ temp1[WIDTH-1:0];
    assign carry = ((in1 ^ in2) ^ in3 ^ in4) & temp1[WIDTH-1:0] | in4 & ~((in1 ^ in2) ^ in3 ^ in4);
    assign cout = temp1[WIDTH];
endmodule




