// Note: The license below is based on the template at:
// http://opensource.org/licenses/BSD-3-Clause
// Copyright (C) 2020 Regents of the University of Texas
//All rights reserved.

// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are
// met:

// o Redistributions of source code must retain the above copyright
//   notice, this list of conditions and the following disclaimer.

// o Redistributions in binary form must reproduce the above copyright
//   notice, this list of conditions and the following disclaimer in the
//   documentation and/or other materials provided with the distribution.

// o Neither the name of the copyright holders nor the names of its
//   contributors may be used to endorse or promote products derived
//   from this software without specific prior written permission.

// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
// A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT
// HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
// SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT
// LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
// DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
// THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

// Original Author(s):
// Mertcan Temel         <mert@utexas.edu>

// DO NOT REMOVE:
// This file is generated by Temel's multiplier generator. Download from https://github.com/temelmertcan/multgen.

// Specification module to help understand what the design implements.
module DT_UB16_KS_16x16_spec (
        input logic [15:0] IN1,
        input logic [15:0] IN2,
        input logic [0:0] IN3, //redundant
        output logic design_is_correct, // is set to 1 iff the output of DT_UB16_KS_16x16 matches its spec.
        output logic [31:0] design_res,
        output logic [31:0] spec_res);
    
    assign spec_res = unsigned'(IN1) * unsigned'(IN2);
    DT_UB16_KS_16x16 mult(IN1, IN2, design_res);
    assign design_is_correct = ((spec_res == design_res) ? 1 : 0);
    
endmodule



module DT_UB16_KS_16x16(
        input logic [15:0] IN1,
        input logic [15:0] IN2,
        output logic [31:0] result);
    
    
// Creating Partial Products 

    wire [16:0] mult = {1'b0, IN1};
    wire [16:0] mcand = {1'b0, IN2};
    wire [19:0] mcand_1x;
    wire [19:0] mcand_2x;
    wire [20:0] mcand_3x;
    wire [19:0] mcand_4x;
    wire [20:0] mcand_5x;
    wire [19:0] mcand_6x;
    wire [20:0] mcand_7x;
    wire [19:0] mcand_8x;
    assign mcand_1x = {{3{mcand[16]}},  mcand};
    assign mcand_2x = {{2{mcand[16]}},  mcand, 1'b0};
    KS_20 calc_mcand_3x (1'b0, mcand_1x, mcand_2x, mcand_3x);
    assign mcand_4x = {{1{mcand[16]}},  mcand, 2'b0};
    KS_20 calc_mcand_5x (1'b0, mcand_1x, mcand_4x, mcand_5x);
    assign mcand_6x = {mcand_3x[18:0], 1'b0};
    KS_20 calc_mcand_7x (1'b1, ~mcand_1x, mcand_8x, mcand_7x);
    assign mcand_8x =  {{0{mcand[16]}},  mcand, 3'b0};
    
    // Booth Radix-16 Partial Products. Multiplier selectors: mult[3] mult[2] mult[1] mult[0] 1'b0
    wire logic select_e_0, select_2x_0, select_3x_0, select_4x_0, select_5x_0, select_6x_0, select_7x_0, select_8x_0, tcomp0, select_ne_0, select_n2x_0, select_n3x_0, select_n4x_0, select_n5x_0, select_n6x_0, select_n7x_0, select_n8x_0, select_0_0;
    assign select_0_0 =  &{mult[3],  mult[2], mult[1], mult[0], 1'b0} | ~|{mult[3],  mult[2], mult[1], mult[0], 1'b0};
    assign select_e_0 = ((~ mult[3]) & (~ mult[2]) & (~ mult[1]) & (mult[0] ^ 1'b0));
    assign select_2x_0 = (~ mult[3]) & (~ mult[2]) & (mult[1] ^ mult[0])& (mult[1] ^ 1'b0);
    assign select_3x_0 = (~ mult[3]) & (~ mult[2]) & mult[1] & (mult[0] ^ 1'b0);
    assign select_4x_0 = (~mult[3]) &  (mult[2] ^ mult[1]) & (mult[2] ^ mult[0])& (mult[2] ^ 1'b0);
    assign select_5x_0 =  (~mult[3]) &  mult[2] & (~mult[1]) & (mult[0] ^ 1'b0);
    assign select_6x_0 = (~mult[3]) & mult[2] & (mult[1] ^ mult[0])& (mult[1] ^ 1'b0);
    assign select_7x_0 =  (~mult[3]) &  mult[2] & mult[1] & (mult[0] ^ 1'b0);
    assign select_8x_0 =  (~mult[3]) &  mult[2] & mult[1] & mult[0] & 1'b0;
    assign select_n8x_0 =  mult[3] &  (~mult[2]) & (~mult[1]) & (~mult[0]) & (~1'b0);
    assign select_n7x_0 = (( mult[3]) & (~ mult[2]) & (~ mult[1]) & (mult[0] ^ 1'b0));
    assign select_n6x_0 = (mult[3]) & (~ mult[2]) & (mult[1] ^ mult[0])& (mult[1] ^ 1'b0);
    assign select_n5x_0 = (mult[3]) & (~ mult[2]) & mult[1] & (mult[0] ^ 1'b0);
    assign select_n4x_0 = (mult[3]) &  (mult[2] ^ mult[1]) & (mult[2] ^ mult[0])& (mult[2] ^ 1'b0);
    assign select_n3x_0 =  (mult[3]) &  mult[2] & (~mult[1]) & (mult[0] ^ 1'b0);
    assign select_n2x_0 = (mult[3]) & mult[2] & (mult[1] ^ mult[0])& (mult[1] ^ 1'b0);
    assign select_ne_0 =  (mult[3]) &  mult[2] & mult[1] & (mult[0] ^ 1'b0);
    reg [19:0] pp_0;
    always @(*) begin
       case (1'b1)
          select_0_0   : pp_0 = 0; 
          select_e_0   : pp_0 = mcand_1x; 
          select_2x_0  : pp_0 = mcand_2x; 
          select_3x_0  : pp_0 = mcand_3x; 
          select_4x_0  : pp_0 = mcand_4x; 
          select_5x_0  : pp_0 = mcand_5x; 
          select_6x_0  : pp_0 = mcand_6x; 
          select_7x_0  : pp_0 = mcand_7x; 
          select_8x_0  : pp_0 = mcand_8x; 
          select_n8x_0 : pp_0 = (~ mcand_8x); 
          select_n7x_0 : pp_0 = (~ mcand_7x); 
          select_n6x_0 : pp_0 = (~ mcand_6x); 
          select_n5x_0 : pp_0 = (~ mcand_5x); 
          select_n4x_0 : pp_0 = (~ mcand_4x); 
          select_n3x_0 : pp_0 = (~ mcand_3x); 
          select_n2x_0 : pp_0 = (~ mcand_2x); 
          select_ne_0  : pp_0 = (~ mcand_1x); 
       endcase 
       pp_0[19] = ~pp_0[19]; // flip the MSB 
    end
    assign tcomp0 = select_ne_0 | select_n8x_0 | select_n7x_0 | select_n6x_0 | select_n5x_0 | select_n4x_0 | select_n3x_0 | select_n2x_0;
    
    // Booth Radix-16 Partial Products. Multiplier selectors: mult[7] mult[6] mult[5] mult[4] mult[3]
    wire logic select_e_1, select_2x_1, select_3x_1, select_4x_1, select_5x_1, select_6x_1, select_7x_1, select_8x_1, tcomp1, select_ne_1, select_n2x_1, select_n3x_1, select_n4x_1, select_n5x_1, select_n6x_1, select_n7x_1, select_n8x_1, select_0_1;
    assign select_0_1 =  &{mult[7],  mult[6], mult[5], mult[4], mult[3]} | ~|{mult[7],  mult[6], mult[5], mult[4], mult[3]};
    assign select_e_1 = ((~ mult[7]) & (~ mult[6]) & (~ mult[5]) & (mult[4] ^ mult[3]));
    assign select_2x_1 = (~ mult[7]) & (~ mult[6]) & (mult[5] ^ mult[4])& (mult[5] ^ mult[3]);
    assign select_3x_1 = (~ mult[7]) & (~ mult[6]) & mult[5] & (mult[4] ^ mult[3]);
    assign select_4x_1 = (~mult[7]) &  (mult[6] ^ mult[5]) & (mult[6] ^ mult[4])& (mult[6] ^ mult[3]);
    assign select_5x_1 =  (~mult[7]) &  mult[6] & (~mult[5]) & (mult[4] ^ mult[3]);
    assign select_6x_1 = (~mult[7]) & mult[6] & (mult[5] ^ mult[4])& (mult[5] ^ mult[3]);
    assign select_7x_1 =  (~mult[7]) &  mult[6] & mult[5] & (mult[4] ^ mult[3]);
    assign select_8x_1 =  (~mult[7]) &  mult[6] & mult[5] & mult[4] & mult[3];
    assign select_n8x_1 =  mult[7] &  (~mult[6]) & (~mult[5]) & (~mult[4]) & (~mult[3]);
    assign select_n7x_1 = (( mult[7]) & (~ mult[6]) & (~ mult[5]) & (mult[4] ^ mult[3]));
    assign select_n6x_1 = (mult[7]) & (~ mult[6]) & (mult[5] ^ mult[4])& (mult[5] ^ mult[3]);
    assign select_n5x_1 = (mult[7]) & (~ mult[6]) & mult[5] & (mult[4] ^ mult[3]);
    assign select_n4x_1 = (mult[7]) &  (mult[6] ^ mult[5]) & (mult[6] ^ mult[4])& (mult[6] ^ mult[3]);
    assign select_n3x_1 =  (mult[7]) &  mult[6] & (~mult[5]) & (mult[4] ^ mult[3]);
    assign select_n2x_1 = (mult[7]) & mult[6] & (mult[5] ^ mult[4])& (mult[5] ^ mult[3]);
    assign select_ne_1 =  (mult[7]) &  mult[6] & mult[5] & (mult[4] ^ mult[3]);
    reg [19:0] pp_1;
    always @(*) begin
       case (1'b1)
          select_0_1   : pp_1 = 0; 
          select_e_1   : pp_1 = mcand_1x; 
          select_2x_1  : pp_1 = mcand_2x; 
          select_3x_1  : pp_1 = mcand_3x; 
          select_4x_1  : pp_1 = mcand_4x; 
          select_5x_1  : pp_1 = mcand_5x; 
          select_6x_1  : pp_1 = mcand_6x; 
          select_7x_1  : pp_1 = mcand_7x; 
          select_8x_1  : pp_1 = mcand_8x; 
          select_n8x_1 : pp_1 = (~ mcand_8x); 
          select_n7x_1 : pp_1 = (~ mcand_7x); 
          select_n6x_1 : pp_1 = (~ mcand_6x); 
          select_n5x_1 : pp_1 = (~ mcand_5x); 
          select_n4x_1 : pp_1 = (~ mcand_4x); 
          select_n3x_1 : pp_1 = (~ mcand_3x); 
          select_n2x_1 : pp_1 = (~ mcand_2x); 
          select_ne_1  : pp_1 = (~ mcand_1x); 
       endcase 
       pp_1[19] = ~pp_1[19]; // flip the MSB 
    end
    assign tcomp1 = select_ne_1 | select_n8x_1 | select_n7x_1 | select_n6x_1 | select_n5x_1 | select_n4x_1 | select_n3x_1 | select_n2x_1;
    
    // Booth Radix-16 Partial Products. Multiplier selectors: mult[11] mult[10] mult[9] mult[8] mult[7]
    wire logic select_e_2, select_2x_2, select_3x_2, select_4x_2, select_5x_2, select_6x_2, select_7x_2, select_8x_2, tcomp2, select_ne_2, select_n2x_2, select_n3x_2, select_n4x_2, select_n5x_2, select_n6x_2, select_n7x_2, select_n8x_2, select_0_2;
    assign select_0_2 =  &{mult[11],  mult[10], mult[9], mult[8], mult[7]} | ~|{mult[11],  mult[10], mult[9], mult[8], mult[7]};
    assign select_e_2 = ((~ mult[11]) & (~ mult[10]) & (~ mult[9]) & (mult[8] ^ mult[7]));
    assign select_2x_2 = (~ mult[11]) & (~ mult[10]) & (mult[9] ^ mult[8])& (mult[9] ^ mult[7]);
    assign select_3x_2 = (~ mult[11]) & (~ mult[10]) & mult[9] & (mult[8] ^ mult[7]);
    assign select_4x_2 = (~mult[11]) &  (mult[10] ^ mult[9]) & (mult[10] ^ mult[8])& (mult[10] ^ mult[7]);
    assign select_5x_2 =  (~mult[11]) &  mult[10] & (~mult[9]) & (mult[8] ^ mult[7]);
    assign select_6x_2 = (~mult[11]) & mult[10] & (mult[9] ^ mult[8])& (mult[9] ^ mult[7]);
    assign select_7x_2 =  (~mult[11]) &  mult[10] & mult[9] & (mult[8] ^ mult[7]);
    assign select_8x_2 =  (~mult[11]) &  mult[10] & mult[9] & mult[8] & mult[7];
    assign select_n8x_2 =  mult[11] &  (~mult[10]) & (~mult[9]) & (~mult[8]) & (~mult[7]);
    assign select_n7x_2 = (( mult[11]) & (~ mult[10]) & (~ mult[9]) & (mult[8] ^ mult[7]));
    assign select_n6x_2 = (mult[11]) & (~ mult[10]) & (mult[9] ^ mult[8])& (mult[9] ^ mult[7]);
    assign select_n5x_2 = (mult[11]) & (~ mult[10]) & mult[9] & (mult[8] ^ mult[7]);
    assign select_n4x_2 = (mult[11]) &  (mult[10] ^ mult[9]) & (mult[10] ^ mult[8])& (mult[10] ^ mult[7]);
    assign select_n3x_2 =  (mult[11]) &  mult[10] & (~mult[9]) & (mult[8] ^ mult[7]);
    assign select_n2x_2 = (mult[11]) & mult[10] & (mult[9] ^ mult[8])& (mult[9] ^ mult[7]);
    assign select_ne_2 =  (mult[11]) &  mult[10] & mult[9] & (mult[8] ^ mult[7]);
    reg [19:0] pp_2;
    always @(*) begin
       case (1'b1)
          select_0_2   : pp_2 = 0; 
          select_e_2   : pp_2 = mcand_1x; 
          select_2x_2  : pp_2 = mcand_2x; 
          select_3x_2  : pp_2 = mcand_3x; 
          select_4x_2  : pp_2 = mcand_4x; 
          select_5x_2  : pp_2 = mcand_5x; 
          select_6x_2  : pp_2 = mcand_6x; 
          select_7x_2  : pp_2 = mcand_7x; 
          select_8x_2  : pp_2 = mcand_8x; 
          select_n8x_2 : pp_2 = (~ mcand_8x); 
          select_n7x_2 : pp_2 = (~ mcand_7x); 
          select_n6x_2 : pp_2 = (~ mcand_6x); 
          select_n5x_2 : pp_2 = (~ mcand_5x); 
          select_n4x_2 : pp_2 = (~ mcand_4x); 
          select_n3x_2 : pp_2 = (~ mcand_3x); 
          select_n2x_2 : pp_2 = (~ mcand_2x); 
          select_ne_2  : pp_2 = (~ mcand_1x); 
       endcase 
       pp_2[19] = ~pp_2[19]; // flip the MSB 
    end
    assign tcomp2 = select_ne_2 | select_n8x_2 | select_n7x_2 | select_n6x_2 | select_n5x_2 | select_n4x_2 | select_n3x_2 | select_n2x_2;
    
    // Booth Radix-16 Partial Products. Multiplier selectors: mult[15] mult[14] mult[13] mult[12] mult[11]
    wire logic select_e_3, select_2x_3, select_3x_3, select_4x_3, select_5x_3, select_6x_3, select_7x_3, select_8x_3, tcomp3, select_ne_3, select_n2x_3, select_n3x_3, select_n4x_3, select_n5x_3, select_n6x_3, select_n7x_3, select_n8x_3, select_0_3;
    assign select_0_3 =  &{mult[15],  mult[14], mult[13], mult[12], mult[11]} | ~|{mult[15],  mult[14], mult[13], mult[12], mult[11]};
    assign select_e_3 = ((~ mult[15]) & (~ mult[14]) & (~ mult[13]) & (mult[12] ^ mult[11]));
    assign select_2x_3 = (~ mult[15]) & (~ mult[14]) & (mult[13] ^ mult[12])& (mult[13] ^ mult[11]);
    assign select_3x_3 = (~ mult[15]) & (~ mult[14]) & mult[13] & (mult[12] ^ mult[11]);
    assign select_4x_3 = (~mult[15]) &  (mult[14] ^ mult[13]) & (mult[14] ^ mult[12])& (mult[14] ^ mult[11]);
    assign select_5x_3 =  (~mult[15]) &  mult[14] & (~mult[13]) & (mult[12] ^ mult[11]);
    assign select_6x_3 = (~mult[15]) & mult[14] & (mult[13] ^ mult[12])& (mult[13] ^ mult[11]);
    assign select_7x_3 =  (~mult[15]) &  mult[14] & mult[13] & (mult[12] ^ mult[11]);
    assign select_8x_3 =  (~mult[15]) &  mult[14] & mult[13] & mult[12] & mult[11];
    assign select_n8x_3 =  mult[15] &  (~mult[14]) & (~mult[13]) & (~mult[12]) & (~mult[11]);
    assign select_n7x_3 = (( mult[15]) & (~ mult[14]) & (~ mult[13]) & (mult[12] ^ mult[11]));
    assign select_n6x_3 = (mult[15]) & (~ mult[14]) & (mult[13] ^ mult[12])& (mult[13] ^ mult[11]);
    assign select_n5x_3 = (mult[15]) & (~ mult[14]) & mult[13] & (mult[12] ^ mult[11]);
    assign select_n4x_3 = (mult[15]) &  (mult[14] ^ mult[13]) & (mult[14] ^ mult[12])& (mult[14] ^ mult[11]);
    assign select_n3x_3 =  (mult[15]) &  mult[14] & (~mult[13]) & (mult[12] ^ mult[11]);
    assign select_n2x_3 = (mult[15]) & mult[14] & (mult[13] ^ mult[12])& (mult[13] ^ mult[11]);
    assign select_ne_3 =  (mult[15]) &  mult[14] & mult[13] & (mult[12] ^ mult[11]);
    reg [19:0] pp_3;
    always @(*) begin
       case (1'b1)
          select_0_3   : pp_3 = 0; 
          select_e_3   : pp_3 = mcand_1x; 
          select_2x_3  : pp_3 = mcand_2x; 
          select_3x_3  : pp_3 = mcand_3x; 
          select_4x_3  : pp_3 = mcand_4x; 
          select_5x_3  : pp_3 = mcand_5x; 
          select_6x_3  : pp_3 = mcand_6x; 
          select_7x_3  : pp_3 = mcand_7x; 
          select_8x_3  : pp_3 = mcand_8x; 
          select_n8x_3 : pp_3 = (~ mcand_8x); 
          select_n7x_3 : pp_3 = (~ mcand_7x); 
          select_n6x_3 : pp_3 = (~ mcand_6x); 
          select_n5x_3 : pp_3 = (~ mcand_5x); 
          select_n4x_3 : pp_3 = (~ mcand_4x); 
          select_n3x_3 : pp_3 = (~ mcand_3x); 
          select_n2x_3 : pp_3 = (~ mcand_2x); 
          select_ne_3  : pp_3 = (~ mcand_1x); 
       endcase 
       pp_3[19] = ~pp_3[19]; // flip the MSB 
    end
    assign tcomp3 = select_ne_3 | select_n8x_3 | select_n7x_3 | select_n6x_3 | select_n5x_3 | select_n4x_3 | select_n3x_3 | select_n2x_3;
    
    // Booth Radix-16 Partial Products. Multiplier selectors: mult[16] mult[16] mult[16] mult[16] mult[15]
    wire logic select_e_4, select_2x_4, select_3x_4, select_4x_4, select_5x_4, select_6x_4, select_7x_4, select_8x_4, tcomp4, select_ne_4, select_n2x_4, select_n3x_4, select_n4x_4, select_n5x_4, select_n6x_4, select_n7x_4, select_n8x_4, select_0_4;
    assign select_0_4 =  &{mult[16],  mult[16], mult[16], mult[16], mult[15]} | ~|{mult[16],  mult[16], mult[16], mult[16], mult[15]};
    assign select_e_4 = ((~ mult[16]) & (~ mult[16]) & (~ mult[16]) & (mult[16] ^ mult[15]));
    assign select_2x_4 = (~ mult[16]) & (~ mult[16]) & (mult[16] ^ mult[16])& (mult[16] ^ mult[15]);
    assign select_3x_4 = (~ mult[16]) & (~ mult[16]) & mult[16] & (mult[16] ^ mult[15]);
    assign select_4x_4 = (~mult[16]) &  (mult[16] ^ mult[16]) & (mult[16] ^ mult[16])& (mult[16] ^ mult[15]);
    assign select_5x_4 =  (~mult[16]) &  mult[16] & (~mult[16]) & (mult[16] ^ mult[15]);
    assign select_6x_4 = (~mult[16]) & mult[16] & (mult[16] ^ mult[16])& (mult[16] ^ mult[15]);
    assign select_7x_4 =  (~mult[16]) &  mult[16] & mult[16] & (mult[16] ^ mult[15]);
    assign select_8x_4 =  (~mult[16]) &  mult[16] & mult[16] & mult[16] & mult[15];
    assign select_n8x_4 =  mult[16] &  (~mult[16]) & (~mult[16]) & (~mult[16]) & (~mult[15]);
    assign select_n7x_4 = (( mult[16]) & (~ mult[16]) & (~ mult[16]) & (mult[16] ^ mult[15]));
    assign select_n6x_4 = (mult[16]) & (~ mult[16]) & (mult[16] ^ mult[16])& (mult[16] ^ mult[15]);
    assign select_n5x_4 = (mult[16]) & (~ mult[16]) & mult[16] & (mult[16] ^ mult[15]);
    assign select_n4x_4 = (mult[16]) &  (mult[16] ^ mult[16]) & (mult[16] ^ mult[16])& (mult[16] ^ mult[15]);
    assign select_n3x_4 =  (mult[16]) &  mult[16] & (~mult[16]) & (mult[16] ^ mult[15]);
    assign select_n2x_4 = (mult[16]) & mult[16] & (mult[16] ^ mult[16])& (mult[16] ^ mult[15]);
    assign select_ne_4 =  (mult[16]) &  mult[16] & mult[16] & (mult[16] ^ mult[15]);
    reg [19:0] pp_4;
    always @(*) begin
       case (1'b1)
          select_0_4   : pp_4 = 0; 
          select_e_4   : pp_4 = mcand_1x; 
          select_2x_4  : pp_4 = mcand_2x; 
          select_3x_4  : pp_4 = mcand_3x; 
          select_4x_4  : pp_4 = mcand_4x; 
          select_5x_4  : pp_4 = mcand_5x; 
          select_6x_4  : pp_4 = mcand_6x; 
          select_7x_4  : pp_4 = mcand_7x; 
          select_8x_4  : pp_4 = mcand_8x; 
          select_n8x_4 : pp_4 = (~ mcand_8x); 
          select_n7x_4 : pp_4 = (~ mcand_7x); 
          select_n6x_4 : pp_4 = (~ mcand_6x); 
          select_n5x_4 : pp_4 = (~ mcand_5x); 
          select_n4x_4 : pp_4 = (~ mcand_4x); 
          select_n3x_4 : pp_4 = (~ mcand_3x); 
          select_n2x_4 : pp_4 = (~ mcand_2x); 
          select_ne_4  : pp_4 = (~ mcand_1x); 
       endcase 
       pp_4[19] = ~pp_4[19]; // flip the MSB 
    end
    assign tcomp4 = select_ne_4 | select_n8x_4 | select_n7x_4 | select_n6x_4 | select_n5x_4 | select_n4x_4 | select_n3x_4 | select_n2x_4;
    
    // The values to be summed in the summation tree, from LSB (left) to MSB:
     // pp_0[0]  pp_0[1]  pp_0[2]  pp_0[3]  pp_0[4]  pp_0[5]  pp_0[6]  pp_0[7]  pp_0[8]  pp_0[9]  pp_0[10] pp_0[11] pp_0[12] pp_0[13] pp_0[14] pp_0[15] pp_0[16] pp_0[17] pp_0[18] pp_0[19]   --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     
     //   --       --       --       --     pp_1[0]  pp_1[1]  pp_1[2]  pp_1[3]  pp_1[4]  pp_1[5]  pp_1[6]  pp_1[7]  pp_1[8]  pp_1[9]  pp_1[10] pp_1[11] pp_1[12] pp_1[13] pp_1[14] pp_1[15] pp_1[16] pp_1[17] pp_1[18] pp_1[19]   --       --       --       --       --       --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --     pp_2[0]  pp_2[1]  pp_2[2]  pp_2[3]  pp_2[4]  pp_2[5]  pp_2[6]  pp_2[7]  pp_2[8]  pp_2[9]  pp_2[10] pp_2[11] pp_2[12] pp_2[13] pp_2[14] pp_2[15] pp_2[16] pp_2[17] pp_2[18] pp_2[19]   --       --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --       --       --       --       --     pp_3[0]  pp_3[1]  pp_3[2]  pp_3[3]  pp_3[4]  pp_3[5]  pp_3[6]  pp_3[7]  pp_3[8]  pp_3[9]  pp_3[10] pp_3[11] pp_3[12] pp_3[13] pp_3[14] pp_3[15] pp_3[16] pp_3[17] pp_3[18] pp_3[19]   --       --       --       --     
     //   --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     pp_4[0]  pp_4[1]  pp_4[2]  pp_4[3]  pp_4[4]  pp_4[5]  pp_4[6]  pp_4[7]  pp_4[8]  pp_4[9]  pp_4[10] pp_4[11] pp_4[12] pp_4[13] pp_4[14] pp_4[15] pp_4[16] pp_4[17] pp_4[18] pp_4[19] 
     // tcomp0     --       --       --     tcomp1     --       --       --     tcomp2     --       --       --     tcomp3     --       --       --     tcomp4     --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     1'b1     1'b1     1'b1     1'b1       --     1'b1     1'b1     1'b1       --     1'b1     1'b1     1'b1       --     1'b1     1'b1     1'b1       --     
    
// Creating Summation Tree 

    
    // Dadda Summation Stage 1
    logic s0 ,c0;
    ha ha0 (pp_0[12], pp_1[8], s0, c0);
    logic s1 ,c1;
    ha ha1 (pp_0[13], pp_1[9], s1, c1);
    logic s2 ,c2;
    ha ha2 (pp_0[14], pp_1[10], s2, c2);
    logic s3 ,c3;
    ha ha3 (pp_0[15], pp_1[11], s3, c3);
    logic s4 ,c4; 
    fa fa4 (pp_0[16], pp_1[12], pp_2[8], s4, c4);
    logic s5 ,c5;
    ha ha5 (pp_3[4], pp_4[0], s5, c5);
    logic s6 ,c6; 
    fa fa6 (pp_0[17], pp_1[13], pp_2[9], s6, c6);
    logic s7 ,c7;
    ha ha7 (pp_3[5], pp_4[1], s7, c7);
    logic s8 ,c8; 
    fa fa8 (pp_0[18], pp_1[14], pp_2[10], s8, c8);
    logic s9 ,c9;
    ha ha9 (pp_3[6], pp_4[2], s9, c9);
    logic s10 ,c10; 
    fa fa10 (pp_0[19], pp_1[15], pp_2[11], s10, c10);
    logic s11 ,c11; 
    fa fa11 (pp_3[7], pp_4[3], 1'b1, s11, c11);
    logic s12 ,c12; 
    fa fa12 (pp_1[16], pp_2[12], pp_3[8], s12, c12);
    logic s13 ,c13;
    ha ha13 (pp_4[4], 1'b1, s13, c13);
    logic s14 ,c14; 
    fa fa14 (pp_1[17], pp_2[13], pp_3[9], s14, c14);
    logic s15 ,c15;
    ha ha15 (pp_4[5], 1'b1, s15, c15);
    logic s16 ,c16; 
    fa fa16 (pp_1[18], pp_2[14], pp_3[10], s16, c16);
    logic s17 ,c17;
    ha ha17 (pp_4[6], 1'b1, s17, c17);
    logic s18 ,c18; 
    fa fa18 (pp_1[19], pp_2[15], pp_3[11], s18, c18);
    logic s19 ,c19;
    ha ha19 (pp_2[16], pp_3[12], s19, c19);
    logic s20 ,c20;
    ha ha20 (pp_2[17], pp_3[13], s20, c20);
    logic s21 ,c21;
    ha ha21 (pp_2[18], pp_3[14], s21, c21);
    
    // Dadda Summation Stage 2
    logic s22 ,c22;
    ha ha22 (pp_0[8], pp_1[4], s22, c22);
    logic s23 ,c23;
    ha ha23 (pp_0[9], pp_1[5], s23, c23);
    logic s24 ,c24;
    ha ha24 (pp_0[10], pp_1[6], s24, c24);
    logic s25 ,c25;
    ha ha25 (pp_0[11], pp_1[7], s25, c25);
    logic s26 ,c26; 
    fa fa26 (pp_2[4], pp_3[0], tcomp3, s26, c26);
    logic s27 ,c27; 
    fa fa27 (pp_2[5], pp_3[1], c0, s27, c27);
    logic s28 ,c28; 
    fa fa28 (pp_2[6], pp_3[2], c1, s28, c28);
    logic s29 ,c29; 
    fa fa29 (pp_2[7], pp_3[3], c2, s29, c29);
    logic s30 ,c30; 
    fa fa30 (tcomp4, c3, s4, s30, c30);
    logic s31 ,c31; 
    fa fa31 (c4, c5, s6, s31, c31);
    logic s32 ,c32; 
    fa fa32 (c6, c7, s8, s32, c32);
    logic s33 ,c33; 
    fa fa33 (c8, c9, s10, s33, c33);
    logic s34 ,c34; 
    fa fa34 (c10, c11, s12, s34, c34);
    logic s35 ,c35; 
    fa fa35 (c12, c13, s14, s35, c35);
    logic s36 ,c36; 
    fa fa36 (c14, c15, s16, s36, c36);
    logic s37 ,c37; 
    fa fa37 (pp_4[7], c16, c17, s37, c37);
    logic s38 ,c38; 
    fa fa38 (pp_4[8], 1'b1, c18, s38, c38);
    logic s39 ,c39; 
    fa fa39 (pp_4[9], 1'b1, c19, s39, c39);
    logic s40 ,c40; 
    fa fa40 (pp_4[10], 1'b1, c20, s40, c40);
    logic s41 ,c41; 
    fa fa41 (pp_2[19], pp_3[15], pp_4[11], s41, c41);
    logic s42 ,c42;
    ha ha42 (pp_3[16], pp_4[12], s42, c42);
    logic s43 ,c43;
    ha ha43 (pp_3[17], pp_4[13], s43, c43);
    logic s44 ,c44;
    ha ha44 (pp_3[18], pp_4[14], s44, c44);
    
    // Dadda Summation Stage 3
    logic s45 ,c45;
    ha ha45 (pp_0[4], pp_1[0], s45, c45);
    logic s46 ,c46;
    ha ha46 (pp_0[5], pp_1[1], s46, c46);
    logic s47 ,c47;
    ha ha47 (pp_0[6], pp_1[2], s47, c47);
    logic s48 ,c48;
    ha ha48 (pp_0[7], pp_1[3], s48, c48);
    logic s49 ,c49; 
    fa fa49 (pp_2[0], tcomp2, s22, s49, c49);
    logic s50 ,c50; 
    fa fa50 (pp_2[1], c22, s23, s50, c50);
    logic s51 ,c51; 
    fa fa51 (pp_2[2], c23, s24, s51, c51);
    logic s52 ,c52; 
    fa fa52 (pp_2[3], c24, s25, s52, c52);
    logic s53 ,c53; 
    fa fa53 (s0, c25, s26, s53, c53);
    logic s54 ,c54; 
    fa fa54 (s1, c26, s27, s54, c54);
    logic s55 ,c55; 
    fa fa55 (s2, c27, s28, s55, c55);
    logic s56 ,c56; 
    fa fa56 (s3, c28, s29, s56, c56);
    logic s57 ,c57; 
    fa fa57 (s5, c29, s30, s57, c57);
    logic s58 ,c58; 
    fa fa58 (s7, c30, s31, s58, c58);
    logic s59 ,c59; 
    fa fa59 (s9, c31, s32, s59, c59);
    logic s60 ,c60; 
    fa fa60 (s11, c32, s33, s60, c60);
    logic s61 ,c61; 
    fa fa61 (s13, c33, s34, s61, c61);
    logic s62 ,c62; 
    fa fa62 (s15, c34, s35, s62, c62);
    logic s63 ,c63; 
    fa fa63 (s17, c35, s36, s63, c63);
    logic s64 ,c64; 
    fa fa64 (s18, c36, s37, s64, c64);
    logic s65 ,c65; 
    fa fa65 (s19, c37, s38, s65, c65);
    logic s66 ,c66; 
    fa fa66 (s20, c38, s39, s66, c66);
    logic s67 ,c67; 
    fa fa67 (s21, c39, s40, s67, c67);
    logic s68 ,c68; 
    fa fa68 (c21, c40, s41, s68, c68);
    logic s69 ,c69; 
    fa fa69 (1'b1, c41, s42, s69, c69);
    logic s70 ,c70; 
    fa fa70 (1'b1, c42, s43, s70, c70);
    logic s71 ,c71; 
    fa fa71 (1'b1, c43, s44, s71, c71);
    logic s72 ,c72; 
    fa fa72 (pp_3[19], pp_4[15], c44, s72, c72);
    
    logic [32:0] adder_result;
    KS_32 final_adder ({c71, c70, c69, c68, c67, c66, c65, c64, c63, c62, c61, c60, c59, c58, c57, c56, c55, c54, c53, c52, c51, c50, c49, c48, c47, c46, c45, tcomp1, pp_0[3], pp_0[2], pp_0[1], pp_0[0] }, {s72, s71, s70, s69, s68, s67, s66, s65, s64, s63, s62, s61, s60, s59, s58, s57, s56, s55, s54, s53, s52, s51, s50, s49, s48, s47, s46, s45, 1'b0, 1'b0, 1'b0, tcomp0 }, adder_result );
    assign result[31:0] = adder_result[31:0];
endmodule



module KS_20 ( 
        input logic carryin,
        input logic [19:0] IN1,
        input logic [19:0] IN2,
        output logic [20:0] OUT);
    
    wire logic [19:0] p_0;
    wire logic [19:0] g_0;
    assign g_0[19:1] = IN1[19:1] & IN2[19:1];
    assign p_0[19:1] = IN1[19:1] ^ IN2[19:1];
    fa m0 (carryin, IN1[0], IN2[0], p_0[0], g_0[0]);
    
// Kogge-Stone Adder 

    
    // KS stage 1
    wire logic p_1_1;
    wire logic g_1_1;
    assign p_1_1 = p_0[1] & p_0[0];
    assign g_1_1 = (p_0[1] & g_0[0]) | g_0[1];
    wire logic p_1_2;
    wire logic g_1_2;
    assign p_1_2 = p_0[2] & p_0[1];
    assign g_1_2 = (p_0[2] & g_0[1]) | g_0[2];
    wire logic p_1_3;
    wire logic g_1_3;
    assign p_1_3 = p_0[3] & p_0[2];
    assign g_1_3 = (p_0[3] & g_0[2]) | g_0[3];
    wire logic p_1_4;
    wire logic g_1_4;
    assign p_1_4 = p_0[4] & p_0[3];
    assign g_1_4 = (p_0[4] & g_0[3]) | g_0[4];
    wire logic p_1_5;
    wire logic g_1_5;
    assign p_1_5 = p_0[5] & p_0[4];
    assign g_1_5 = (p_0[5] & g_0[4]) | g_0[5];
    wire logic p_1_6;
    wire logic g_1_6;
    assign p_1_6 = p_0[6] & p_0[5];
    assign g_1_6 = (p_0[6] & g_0[5]) | g_0[6];
    wire logic p_1_7;
    wire logic g_1_7;
    assign p_1_7 = p_0[7] & p_0[6];
    assign g_1_7 = (p_0[7] & g_0[6]) | g_0[7];
    wire logic p_1_8;
    wire logic g_1_8;
    assign p_1_8 = p_0[8] & p_0[7];
    assign g_1_8 = (p_0[8] & g_0[7]) | g_0[8];
    wire logic p_1_9;
    wire logic g_1_9;
    assign p_1_9 = p_0[9] & p_0[8];
    assign g_1_9 = (p_0[9] & g_0[8]) | g_0[9];
    wire logic p_1_10;
    wire logic g_1_10;
    assign p_1_10 = p_0[10] & p_0[9];
    assign g_1_10 = (p_0[10] & g_0[9]) | g_0[10];
    wire logic p_1_11;
    wire logic g_1_11;
    assign p_1_11 = p_0[11] & p_0[10];
    assign g_1_11 = (p_0[11] & g_0[10]) | g_0[11];
    wire logic p_1_12;
    wire logic g_1_12;
    assign p_1_12 = p_0[12] & p_0[11];
    assign g_1_12 = (p_0[12] & g_0[11]) | g_0[12];
    wire logic p_1_13;
    wire logic g_1_13;
    assign p_1_13 = p_0[13] & p_0[12];
    assign g_1_13 = (p_0[13] & g_0[12]) | g_0[13];
    wire logic p_1_14;
    wire logic g_1_14;
    assign p_1_14 = p_0[14] & p_0[13];
    assign g_1_14 = (p_0[14] & g_0[13]) | g_0[14];
    wire logic p_1_15;
    wire logic g_1_15;
    assign p_1_15 = p_0[15] & p_0[14];
    assign g_1_15 = (p_0[15] & g_0[14]) | g_0[15];
    wire logic p_1_16;
    wire logic g_1_16;
    assign p_1_16 = p_0[16] & p_0[15];
    assign g_1_16 = (p_0[16] & g_0[15]) | g_0[16];
    wire logic p_1_17;
    wire logic g_1_17;
    assign p_1_17 = p_0[17] & p_0[16];
    assign g_1_17 = (p_0[17] & g_0[16]) | g_0[17];
    wire logic p_1_18;
    wire logic g_1_18;
    assign p_1_18 = p_0[18] & p_0[17];
    assign g_1_18 = (p_0[18] & g_0[17]) | g_0[18];
    wire logic p_1_19;
    wire logic g_1_19;
    assign p_1_19 = p_0[19] & p_0[18];
    assign g_1_19 = (p_0[19] & g_0[18]) | g_0[19];
    
    // KS stage 2
    wire logic p_2_2;
    wire logic g_2_2;
    assign p_2_2 = p_1_2 & p_0[0];
    assign g_2_2 = (p_1_2 & g_0[0]) | g_1_2;
    wire logic p_2_3;
    wire logic g_2_3;
    assign p_2_3 = p_1_3 & p_1_1;
    assign g_2_3 = (p_1_3 & g_1_1) | g_1_3;
    wire logic p_2_4;
    wire logic g_2_4;
    assign p_2_4 = p_1_4 & p_1_2;
    assign g_2_4 = (p_1_4 & g_1_2) | g_1_4;
    wire logic p_2_5;
    wire logic g_2_5;
    assign p_2_5 = p_1_5 & p_1_3;
    assign g_2_5 = (p_1_5 & g_1_3) | g_1_5;
    wire logic p_2_6;
    wire logic g_2_6;
    assign p_2_6 = p_1_6 & p_1_4;
    assign g_2_6 = (p_1_6 & g_1_4) | g_1_6;
    wire logic p_2_7;
    wire logic g_2_7;
    assign p_2_7 = p_1_7 & p_1_5;
    assign g_2_7 = (p_1_7 & g_1_5) | g_1_7;
    wire logic p_2_8;
    wire logic g_2_8;
    assign p_2_8 = p_1_8 & p_1_6;
    assign g_2_8 = (p_1_8 & g_1_6) | g_1_8;
    wire logic p_2_9;
    wire logic g_2_9;
    assign p_2_9 = p_1_9 & p_1_7;
    assign g_2_9 = (p_1_9 & g_1_7) | g_1_9;
    wire logic p_2_10;
    wire logic g_2_10;
    assign p_2_10 = p_1_10 & p_1_8;
    assign g_2_10 = (p_1_10 & g_1_8) | g_1_10;
    wire logic p_2_11;
    wire logic g_2_11;
    assign p_2_11 = p_1_11 & p_1_9;
    assign g_2_11 = (p_1_11 & g_1_9) | g_1_11;
    wire logic p_2_12;
    wire logic g_2_12;
    assign p_2_12 = p_1_12 & p_1_10;
    assign g_2_12 = (p_1_12 & g_1_10) | g_1_12;
    wire logic p_2_13;
    wire logic g_2_13;
    assign p_2_13 = p_1_13 & p_1_11;
    assign g_2_13 = (p_1_13 & g_1_11) | g_1_13;
    wire logic p_2_14;
    wire logic g_2_14;
    assign p_2_14 = p_1_14 & p_1_12;
    assign g_2_14 = (p_1_14 & g_1_12) | g_1_14;
    wire logic p_2_15;
    wire logic g_2_15;
    assign p_2_15 = p_1_15 & p_1_13;
    assign g_2_15 = (p_1_15 & g_1_13) | g_1_15;
    wire logic p_2_16;
    wire logic g_2_16;
    assign p_2_16 = p_1_16 & p_1_14;
    assign g_2_16 = (p_1_16 & g_1_14) | g_1_16;
    wire logic p_2_17;
    wire logic g_2_17;
    assign p_2_17 = p_1_17 & p_1_15;
    assign g_2_17 = (p_1_17 & g_1_15) | g_1_17;
    wire logic p_2_18;
    wire logic g_2_18;
    assign p_2_18 = p_1_18 & p_1_16;
    assign g_2_18 = (p_1_18 & g_1_16) | g_1_18;
    wire logic p_2_19;
    wire logic g_2_19;
    assign p_2_19 = p_1_19 & p_1_17;
    assign g_2_19 = (p_1_19 & g_1_17) | g_1_19;
    
    // KS stage 3
    wire logic p_3_4;
    wire logic g_3_4;
    assign p_3_4 = p_2_4 & p_0[0];
    assign g_3_4 = (p_2_4 & g_0[0]) | g_2_4;
    wire logic p_3_5;
    wire logic g_3_5;
    assign p_3_5 = p_2_5 & p_1_1;
    assign g_3_5 = (p_2_5 & g_1_1) | g_2_5;
    wire logic p_3_6;
    wire logic g_3_6;
    assign p_3_6 = p_2_6 & p_2_2;
    assign g_3_6 = (p_2_6 & g_2_2) | g_2_6;
    wire logic p_3_7;
    wire logic g_3_7;
    assign p_3_7 = p_2_7 & p_2_3;
    assign g_3_7 = (p_2_7 & g_2_3) | g_2_7;
    wire logic p_3_8;
    wire logic g_3_8;
    assign p_3_8 = p_2_8 & p_2_4;
    assign g_3_8 = (p_2_8 & g_2_4) | g_2_8;
    wire logic p_3_9;
    wire logic g_3_9;
    assign p_3_9 = p_2_9 & p_2_5;
    assign g_3_9 = (p_2_9 & g_2_5) | g_2_9;
    wire logic p_3_10;
    wire logic g_3_10;
    assign p_3_10 = p_2_10 & p_2_6;
    assign g_3_10 = (p_2_10 & g_2_6) | g_2_10;
    wire logic p_3_11;
    wire logic g_3_11;
    assign p_3_11 = p_2_11 & p_2_7;
    assign g_3_11 = (p_2_11 & g_2_7) | g_2_11;
    wire logic p_3_12;
    wire logic g_3_12;
    assign p_3_12 = p_2_12 & p_2_8;
    assign g_3_12 = (p_2_12 & g_2_8) | g_2_12;
    wire logic p_3_13;
    wire logic g_3_13;
    assign p_3_13 = p_2_13 & p_2_9;
    assign g_3_13 = (p_2_13 & g_2_9) | g_2_13;
    wire logic p_3_14;
    wire logic g_3_14;
    assign p_3_14 = p_2_14 & p_2_10;
    assign g_3_14 = (p_2_14 & g_2_10) | g_2_14;
    wire logic p_3_15;
    wire logic g_3_15;
    assign p_3_15 = p_2_15 & p_2_11;
    assign g_3_15 = (p_2_15 & g_2_11) | g_2_15;
    wire logic p_3_16;
    wire logic g_3_16;
    assign p_3_16 = p_2_16 & p_2_12;
    assign g_3_16 = (p_2_16 & g_2_12) | g_2_16;
    wire logic p_3_17;
    wire logic g_3_17;
    assign p_3_17 = p_2_17 & p_2_13;
    assign g_3_17 = (p_2_17 & g_2_13) | g_2_17;
    wire logic p_3_18;
    wire logic g_3_18;
    assign p_3_18 = p_2_18 & p_2_14;
    assign g_3_18 = (p_2_18 & g_2_14) | g_2_18;
    wire logic p_3_19;
    wire logic g_3_19;
    assign p_3_19 = p_2_19 & p_2_15;
    assign g_3_19 = (p_2_19 & g_2_15) | g_2_19;
    
    // KS stage 4
    wire logic p_4_8;
    wire logic g_4_8;
    assign p_4_8 = p_3_8 & p_0[0];
    assign g_4_8 = (p_3_8 & g_0[0]) | g_3_8;
    wire logic p_4_9;
    wire logic g_4_9;
    assign p_4_9 = p_3_9 & p_1_1;
    assign g_4_9 = (p_3_9 & g_1_1) | g_3_9;
    wire logic p_4_10;
    wire logic g_4_10;
    assign p_4_10 = p_3_10 & p_2_2;
    assign g_4_10 = (p_3_10 & g_2_2) | g_3_10;
    wire logic p_4_11;
    wire logic g_4_11;
    assign p_4_11 = p_3_11 & p_2_3;
    assign g_4_11 = (p_3_11 & g_2_3) | g_3_11;
    wire logic p_4_12;
    wire logic g_4_12;
    assign p_4_12 = p_3_12 & p_3_4;
    assign g_4_12 = (p_3_12 & g_3_4) | g_3_12;
    wire logic p_4_13;
    wire logic g_4_13;
    assign p_4_13 = p_3_13 & p_3_5;
    assign g_4_13 = (p_3_13 & g_3_5) | g_3_13;
    wire logic p_4_14;
    wire logic g_4_14;
    assign p_4_14 = p_3_14 & p_3_6;
    assign g_4_14 = (p_3_14 & g_3_6) | g_3_14;
    wire logic p_4_15;
    wire logic g_4_15;
    assign p_4_15 = p_3_15 & p_3_7;
    assign g_4_15 = (p_3_15 & g_3_7) | g_3_15;
    wire logic p_4_16;
    wire logic g_4_16;
    assign p_4_16 = p_3_16 & p_3_8;
    assign g_4_16 = (p_3_16 & g_3_8) | g_3_16;
    wire logic p_4_17;
    wire logic g_4_17;
    assign p_4_17 = p_3_17 & p_3_9;
    assign g_4_17 = (p_3_17 & g_3_9) | g_3_17;
    wire logic p_4_18;
    wire logic g_4_18;
    assign p_4_18 = p_3_18 & p_3_10;
    assign g_4_18 = (p_3_18 & g_3_10) | g_3_18;
    wire logic p_4_19;
    wire logic g_4_19;
    assign p_4_19 = p_3_19 & p_3_11;
    assign g_4_19 = (p_3_19 & g_3_11) | g_3_19;
    
    // KS stage 5
    wire logic p_5_16;
    wire logic g_5_16;
    assign p_5_16 = p_4_16 & p_0[0];
    assign g_5_16 = (p_4_16 & g_0[0]) | g_4_16;
    wire logic p_5_17;
    wire logic g_5_17;
    assign p_5_17 = p_4_17 & p_1_1;
    assign g_5_17 = (p_4_17 & g_1_1) | g_4_17;
    wire logic p_5_18;
    wire logic g_5_18;
    assign p_5_18 = p_4_18 & p_2_2;
    assign g_5_18 = (p_4_18 & g_2_2) | g_4_18;
    wire logic p_5_19;
    wire logic g_5_19;
    assign p_5_19 = p_4_19 & p_2_3;
    assign g_5_19 = (p_4_19 & g_2_3) | g_4_19;
    
    // KS postprocess 
    assign OUT[0] = p_0[0];
    assign OUT[1] = p_0[1] ^ g_0[0];
    assign OUT[2] = p_0[2] ^ g_1_1;
    assign OUT[3] = p_0[3] ^ g_2_2;
    assign OUT[4] = p_0[4] ^ g_2_3;
    assign OUT[5] = p_0[5] ^ g_3_4;
    assign OUT[6] = p_0[6] ^ g_3_5;
    assign OUT[7] = p_0[7] ^ g_3_6;
    assign OUT[8] = p_0[8] ^ g_3_7;
    assign OUT[9] = p_0[9] ^ g_4_8;
    assign OUT[10] = p_0[10] ^ g_4_9;
    assign OUT[11] = p_0[11] ^ g_4_10;
    assign OUT[12] = p_0[12] ^ g_4_11;
    assign OUT[13] = p_0[13] ^ g_4_12;
    assign OUT[14] = p_0[14] ^ g_4_13;
    assign OUT[15] = p_0[15] ^ g_4_14;
    assign OUT[16] = p_0[16] ^ g_4_15;
    assign OUT[17] = p_0[17] ^ g_5_16;
    assign OUT[18] = p_0[18] ^ g_5_17;
    assign OUT[19] = p_0[19] ^ g_5_18;
    assign OUT[20] = g_5_19;
endmodule

module KS_20_spec (
        input logic carryin,
        input logic [19:0] IN1,
        input logic [19:0] IN2,
        output logic adder_correct,
        output logic [20:0] spec_res);
    
    assign spec_res = IN1 + IN2 + carryin;
    wire [20:0] adder_res;
    KS_20 adder(carryin, IN1, IN2, adder_res);
    assign adder_correct = ((spec_res == adder_res) ? 1 : 0);
    
endmodule



module KS_32 ( 
        input logic [31:0] IN1,
        input logic [31:0] IN2,
        output logic [32:0] OUT);
    
    wire logic [31:0] p_0;
    wire logic [31:0] g_0;
    assign g_0 = IN1 & IN2;
    assign p_0 = IN1 ^ IN2;
    
// Kogge-Stone Adder 

    
    // KS stage 1
    wire logic p_1_1;
    wire logic g_1_1;
    assign p_1_1 = p_0[1] & p_0[0];
    assign g_1_1 = (p_0[1] & g_0[0]) | g_0[1];
    wire logic p_1_2;
    wire logic g_1_2;
    assign p_1_2 = p_0[2] & p_0[1];
    assign g_1_2 = (p_0[2] & g_0[1]) | g_0[2];
    wire logic p_1_3;
    wire logic g_1_3;
    assign p_1_3 = p_0[3] & p_0[2];
    assign g_1_3 = (p_0[3] & g_0[2]) | g_0[3];
    wire logic p_1_4;
    wire logic g_1_4;
    assign p_1_4 = p_0[4] & p_0[3];
    assign g_1_4 = (p_0[4] & g_0[3]) | g_0[4];
    wire logic p_1_5;
    wire logic g_1_5;
    assign p_1_5 = p_0[5] & p_0[4];
    assign g_1_5 = (p_0[5] & g_0[4]) | g_0[5];
    wire logic p_1_6;
    wire logic g_1_6;
    assign p_1_6 = p_0[6] & p_0[5];
    assign g_1_6 = (p_0[6] & g_0[5]) | g_0[6];
    wire logic p_1_7;
    wire logic g_1_7;
    assign p_1_7 = p_0[7] & p_0[6];
    assign g_1_7 = (p_0[7] & g_0[6]) | g_0[7];
    wire logic p_1_8;
    wire logic g_1_8;
    assign p_1_8 = p_0[8] & p_0[7];
    assign g_1_8 = (p_0[8] & g_0[7]) | g_0[8];
    wire logic p_1_9;
    wire logic g_1_9;
    assign p_1_9 = p_0[9] & p_0[8];
    assign g_1_9 = (p_0[9] & g_0[8]) | g_0[9];
    wire logic p_1_10;
    wire logic g_1_10;
    assign p_1_10 = p_0[10] & p_0[9];
    assign g_1_10 = (p_0[10] & g_0[9]) | g_0[10];
    wire logic p_1_11;
    wire logic g_1_11;
    assign p_1_11 = p_0[11] & p_0[10];
    assign g_1_11 = (p_0[11] & g_0[10]) | g_0[11];
    wire logic p_1_12;
    wire logic g_1_12;
    assign p_1_12 = p_0[12] & p_0[11];
    assign g_1_12 = (p_0[12] & g_0[11]) | g_0[12];
    wire logic p_1_13;
    wire logic g_1_13;
    assign p_1_13 = p_0[13] & p_0[12];
    assign g_1_13 = (p_0[13] & g_0[12]) | g_0[13];
    wire logic p_1_14;
    wire logic g_1_14;
    assign p_1_14 = p_0[14] & p_0[13];
    assign g_1_14 = (p_0[14] & g_0[13]) | g_0[14];
    wire logic p_1_15;
    wire logic g_1_15;
    assign p_1_15 = p_0[15] & p_0[14];
    assign g_1_15 = (p_0[15] & g_0[14]) | g_0[15];
    wire logic p_1_16;
    wire logic g_1_16;
    assign p_1_16 = p_0[16] & p_0[15];
    assign g_1_16 = (p_0[16] & g_0[15]) | g_0[16];
    wire logic p_1_17;
    wire logic g_1_17;
    assign p_1_17 = p_0[17] & p_0[16];
    assign g_1_17 = (p_0[17] & g_0[16]) | g_0[17];
    wire logic p_1_18;
    wire logic g_1_18;
    assign p_1_18 = p_0[18] & p_0[17];
    assign g_1_18 = (p_0[18] & g_0[17]) | g_0[18];
    wire logic p_1_19;
    wire logic g_1_19;
    assign p_1_19 = p_0[19] & p_0[18];
    assign g_1_19 = (p_0[19] & g_0[18]) | g_0[19];
    wire logic p_1_20;
    wire logic g_1_20;
    assign p_1_20 = p_0[20] & p_0[19];
    assign g_1_20 = (p_0[20] & g_0[19]) | g_0[20];
    wire logic p_1_21;
    wire logic g_1_21;
    assign p_1_21 = p_0[21] & p_0[20];
    assign g_1_21 = (p_0[21] & g_0[20]) | g_0[21];
    wire logic p_1_22;
    wire logic g_1_22;
    assign p_1_22 = p_0[22] & p_0[21];
    assign g_1_22 = (p_0[22] & g_0[21]) | g_0[22];
    wire logic p_1_23;
    wire logic g_1_23;
    assign p_1_23 = p_0[23] & p_0[22];
    assign g_1_23 = (p_0[23] & g_0[22]) | g_0[23];
    wire logic p_1_24;
    wire logic g_1_24;
    assign p_1_24 = p_0[24] & p_0[23];
    assign g_1_24 = (p_0[24] & g_0[23]) | g_0[24];
    wire logic p_1_25;
    wire logic g_1_25;
    assign p_1_25 = p_0[25] & p_0[24];
    assign g_1_25 = (p_0[25] & g_0[24]) | g_0[25];
    wire logic p_1_26;
    wire logic g_1_26;
    assign p_1_26 = p_0[26] & p_0[25];
    assign g_1_26 = (p_0[26] & g_0[25]) | g_0[26];
    wire logic p_1_27;
    wire logic g_1_27;
    assign p_1_27 = p_0[27] & p_0[26];
    assign g_1_27 = (p_0[27] & g_0[26]) | g_0[27];
    wire logic p_1_28;
    wire logic g_1_28;
    assign p_1_28 = p_0[28] & p_0[27];
    assign g_1_28 = (p_0[28] & g_0[27]) | g_0[28];
    wire logic p_1_29;
    wire logic g_1_29;
    assign p_1_29 = p_0[29] & p_0[28];
    assign g_1_29 = (p_0[29] & g_0[28]) | g_0[29];
    wire logic p_1_30;
    wire logic g_1_30;
    assign p_1_30 = p_0[30] & p_0[29];
    assign g_1_30 = (p_0[30] & g_0[29]) | g_0[30];
    wire logic p_1_31;
    wire logic g_1_31;
    assign p_1_31 = p_0[31] & p_0[30];
    assign g_1_31 = (p_0[31] & g_0[30]) | g_0[31];
    
    // KS stage 2
    wire logic p_2_2;
    wire logic g_2_2;
    assign p_2_2 = p_1_2 & p_0[0];
    assign g_2_2 = (p_1_2 & g_0[0]) | g_1_2;
    wire logic p_2_3;
    wire logic g_2_3;
    assign p_2_3 = p_1_3 & p_1_1;
    assign g_2_3 = (p_1_3 & g_1_1) | g_1_3;
    wire logic p_2_4;
    wire logic g_2_4;
    assign p_2_4 = p_1_4 & p_1_2;
    assign g_2_4 = (p_1_4 & g_1_2) | g_1_4;
    wire logic p_2_5;
    wire logic g_2_5;
    assign p_2_5 = p_1_5 & p_1_3;
    assign g_2_5 = (p_1_5 & g_1_3) | g_1_5;
    wire logic p_2_6;
    wire logic g_2_6;
    assign p_2_6 = p_1_6 & p_1_4;
    assign g_2_6 = (p_1_6 & g_1_4) | g_1_6;
    wire logic p_2_7;
    wire logic g_2_7;
    assign p_2_7 = p_1_7 & p_1_5;
    assign g_2_7 = (p_1_7 & g_1_5) | g_1_7;
    wire logic p_2_8;
    wire logic g_2_8;
    assign p_2_8 = p_1_8 & p_1_6;
    assign g_2_8 = (p_1_8 & g_1_6) | g_1_8;
    wire logic p_2_9;
    wire logic g_2_9;
    assign p_2_9 = p_1_9 & p_1_7;
    assign g_2_9 = (p_1_9 & g_1_7) | g_1_9;
    wire logic p_2_10;
    wire logic g_2_10;
    assign p_2_10 = p_1_10 & p_1_8;
    assign g_2_10 = (p_1_10 & g_1_8) | g_1_10;
    wire logic p_2_11;
    wire logic g_2_11;
    assign p_2_11 = p_1_11 & p_1_9;
    assign g_2_11 = (p_1_11 & g_1_9) | g_1_11;
    wire logic p_2_12;
    wire logic g_2_12;
    assign p_2_12 = p_1_12 & p_1_10;
    assign g_2_12 = (p_1_12 & g_1_10) | g_1_12;
    wire logic p_2_13;
    wire logic g_2_13;
    assign p_2_13 = p_1_13 & p_1_11;
    assign g_2_13 = (p_1_13 & g_1_11) | g_1_13;
    wire logic p_2_14;
    wire logic g_2_14;
    assign p_2_14 = p_1_14 & p_1_12;
    assign g_2_14 = (p_1_14 & g_1_12) | g_1_14;
    wire logic p_2_15;
    wire logic g_2_15;
    assign p_2_15 = p_1_15 & p_1_13;
    assign g_2_15 = (p_1_15 & g_1_13) | g_1_15;
    wire logic p_2_16;
    wire logic g_2_16;
    assign p_2_16 = p_1_16 & p_1_14;
    assign g_2_16 = (p_1_16 & g_1_14) | g_1_16;
    wire logic p_2_17;
    wire logic g_2_17;
    assign p_2_17 = p_1_17 & p_1_15;
    assign g_2_17 = (p_1_17 & g_1_15) | g_1_17;
    wire logic p_2_18;
    wire logic g_2_18;
    assign p_2_18 = p_1_18 & p_1_16;
    assign g_2_18 = (p_1_18 & g_1_16) | g_1_18;
    wire logic p_2_19;
    wire logic g_2_19;
    assign p_2_19 = p_1_19 & p_1_17;
    assign g_2_19 = (p_1_19 & g_1_17) | g_1_19;
    wire logic p_2_20;
    wire logic g_2_20;
    assign p_2_20 = p_1_20 & p_1_18;
    assign g_2_20 = (p_1_20 & g_1_18) | g_1_20;
    wire logic p_2_21;
    wire logic g_2_21;
    assign p_2_21 = p_1_21 & p_1_19;
    assign g_2_21 = (p_1_21 & g_1_19) | g_1_21;
    wire logic p_2_22;
    wire logic g_2_22;
    assign p_2_22 = p_1_22 & p_1_20;
    assign g_2_22 = (p_1_22 & g_1_20) | g_1_22;
    wire logic p_2_23;
    wire logic g_2_23;
    assign p_2_23 = p_1_23 & p_1_21;
    assign g_2_23 = (p_1_23 & g_1_21) | g_1_23;
    wire logic p_2_24;
    wire logic g_2_24;
    assign p_2_24 = p_1_24 & p_1_22;
    assign g_2_24 = (p_1_24 & g_1_22) | g_1_24;
    wire logic p_2_25;
    wire logic g_2_25;
    assign p_2_25 = p_1_25 & p_1_23;
    assign g_2_25 = (p_1_25 & g_1_23) | g_1_25;
    wire logic p_2_26;
    wire logic g_2_26;
    assign p_2_26 = p_1_26 & p_1_24;
    assign g_2_26 = (p_1_26 & g_1_24) | g_1_26;
    wire logic p_2_27;
    wire logic g_2_27;
    assign p_2_27 = p_1_27 & p_1_25;
    assign g_2_27 = (p_1_27 & g_1_25) | g_1_27;
    wire logic p_2_28;
    wire logic g_2_28;
    assign p_2_28 = p_1_28 & p_1_26;
    assign g_2_28 = (p_1_28 & g_1_26) | g_1_28;
    wire logic p_2_29;
    wire logic g_2_29;
    assign p_2_29 = p_1_29 & p_1_27;
    assign g_2_29 = (p_1_29 & g_1_27) | g_1_29;
    wire logic p_2_30;
    wire logic g_2_30;
    assign p_2_30 = p_1_30 & p_1_28;
    assign g_2_30 = (p_1_30 & g_1_28) | g_1_30;
    wire logic p_2_31;
    wire logic g_2_31;
    assign p_2_31 = p_1_31 & p_1_29;
    assign g_2_31 = (p_1_31 & g_1_29) | g_1_31;
    
    // KS stage 3
    wire logic p_3_4;
    wire logic g_3_4;
    assign p_3_4 = p_2_4 & p_0[0];
    assign g_3_4 = (p_2_4 & g_0[0]) | g_2_4;
    wire logic p_3_5;
    wire logic g_3_5;
    assign p_3_5 = p_2_5 & p_1_1;
    assign g_3_5 = (p_2_5 & g_1_1) | g_2_5;
    wire logic p_3_6;
    wire logic g_3_6;
    assign p_3_6 = p_2_6 & p_2_2;
    assign g_3_6 = (p_2_6 & g_2_2) | g_2_6;
    wire logic p_3_7;
    wire logic g_3_7;
    assign p_3_7 = p_2_7 & p_2_3;
    assign g_3_7 = (p_2_7 & g_2_3) | g_2_7;
    wire logic p_3_8;
    wire logic g_3_8;
    assign p_3_8 = p_2_8 & p_2_4;
    assign g_3_8 = (p_2_8 & g_2_4) | g_2_8;
    wire logic p_3_9;
    wire logic g_3_9;
    assign p_3_9 = p_2_9 & p_2_5;
    assign g_3_9 = (p_2_9 & g_2_5) | g_2_9;
    wire logic p_3_10;
    wire logic g_3_10;
    assign p_3_10 = p_2_10 & p_2_6;
    assign g_3_10 = (p_2_10 & g_2_6) | g_2_10;
    wire logic p_3_11;
    wire logic g_3_11;
    assign p_3_11 = p_2_11 & p_2_7;
    assign g_3_11 = (p_2_11 & g_2_7) | g_2_11;
    wire logic p_3_12;
    wire logic g_3_12;
    assign p_3_12 = p_2_12 & p_2_8;
    assign g_3_12 = (p_2_12 & g_2_8) | g_2_12;
    wire logic p_3_13;
    wire logic g_3_13;
    assign p_3_13 = p_2_13 & p_2_9;
    assign g_3_13 = (p_2_13 & g_2_9) | g_2_13;
    wire logic p_3_14;
    wire logic g_3_14;
    assign p_3_14 = p_2_14 & p_2_10;
    assign g_3_14 = (p_2_14 & g_2_10) | g_2_14;
    wire logic p_3_15;
    wire logic g_3_15;
    assign p_3_15 = p_2_15 & p_2_11;
    assign g_3_15 = (p_2_15 & g_2_11) | g_2_15;
    wire logic p_3_16;
    wire logic g_3_16;
    assign p_3_16 = p_2_16 & p_2_12;
    assign g_3_16 = (p_2_16 & g_2_12) | g_2_16;
    wire logic p_3_17;
    wire logic g_3_17;
    assign p_3_17 = p_2_17 & p_2_13;
    assign g_3_17 = (p_2_17 & g_2_13) | g_2_17;
    wire logic p_3_18;
    wire logic g_3_18;
    assign p_3_18 = p_2_18 & p_2_14;
    assign g_3_18 = (p_2_18 & g_2_14) | g_2_18;
    wire logic p_3_19;
    wire logic g_3_19;
    assign p_3_19 = p_2_19 & p_2_15;
    assign g_3_19 = (p_2_19 & g_2_15) | g_2_19;
    wire logic p_3_20;
    wire logic g_3_20;
    assign p_3_20 = p_2_20 & p_2_16;
    assign g_3_20 = (p_2_20 & g_2_16) | g_2_20;
    wire logic p_3_21;
    wire logic g_3_21;
    assign p_3_21 = p_2_21 & p_2_17;
    assign g_3_21 = (p_2_21 & g_2_17) | g_2_21;
    wire logic p_3_22;
    wire logic g_3_22;
    assign p_3_22 = p_2_22 & p_2_18;
    assign g_3_22 = (p_2_22 & g_2_18) | g_2_22;
    wire logic p_3_23;
    wire logic g_3_23;
    assign p_3_23 = p_2_23 & p_2_19;
    assign g_3_23 = (p_2_23 & g_2_19) | g_2_23;
    wire logic p_3_24;
    wire logic g_3_24;
    assign p_3_24 = p_2_24 & p_2_20;
    assign g_3_24 = (p_2_24 & g_2_20) | g_2_24;
    wire logic p_3_25;
    wire logic g_3_25;
    assign p_3_25 = p_2_25 & p_2_21;
    assign g_3_25 = (p_2_25 & g_2_21) | g_2_25;
    wire logic p_3_26;
    wire logic g_3_26;
    assign p_3_26 = p_2_26 & p_2_22;
    assign g_3_26 = (p_2_26 & g_2_22) | g_2_26;
    wire logic p_3_27;
    wire logic g_3_27;
    assign p_3_27 = p_2_27 & p_2_23;
    assign g_3_27 = (p_2_27 & g_2_23) | g_2_27;
    wire logic p_3_28;
    wire logic g_3_28;
    assign p_3_28 = p_2_28 & p_2_24;
    assign g_3_28 = (p_2_28 & g_2_24) | g_2_28;
    wire logic p_3_29;
    wire logic g_3_29;
    assign p_3_29 = p_2_29 & p_2_25;
    assign g_3_29 = (p_2_29 & g_2_25) | g_2_29;
    wire logic p_3_30;
    wire logic g_3_30;
    assign p_3_30 = p_2_30 & p_2_26;
    assign g_3_30 = (p_2_30 & g_2_26) | g_2_30;
    wire logic p_3_31;
    wire logic g_3_31;
    assign p_3_31 = p_2_31 & p_2_27;
    assign g_3_31 = (p_2_31 & g_2_27) | g_2_31;
    
    // KS stage 4
    wire logic p_4_8;
    wire logic g_4_8;
    assign p_4_8 = p_3_8 & p_0[0];
    assign g_4_8 = (p_3_8 & g_0[0]) | g_3_8;
    wire logic p_4_9;
    wire logic g_4_9;
    assign p_4_9 = p_3_9 & p_1_1;
    assign g_4_9 = (p_3_9 & g_1_1) | g_3_9;
    wire logic p_4_10;
    wire logic g_4_10;
    assign p_4_10 = p_3_10 & p_2_2;
    assign g_4_10 = (p_3_10 & g_2_2) | g_3_10;
    wire logic p_4_11;
    wire logic g_4_11;
    assign p_4_11 = p_3_11 & p_2_3;
    assign g_4_11 = (p_3_11 & g_2_3) | g_3_11;
    wire logic p_4_12;
    wire logic g_4_12;
    assign p_4_12 = p_3_12 & p_3_4;
    assign g_4_12 = (p_3_12 & g_3_4) | g_3_12;
    wire logic p_4_13;
    wire logic g_4_13;
    assign p_4_13 = p_3_13 & p_3_5;
    assign g_4_13 = (p_3_13 & g_3_5) | g_3_13;
    wire logic p_4_14;
    wire logic g_4_14;
    assign p_4_14 = p_3_14 & p_3_6;
    assign g_4_14 = (p_3_14 & g_3_6) | g_3_14;
    wire logic p_4_15;
    wire logic g_4_15;
    assign p_4_15 = p_3_15 & p_3_7;
    assign g_4_15 = (p_3_15 & g_3_7) | g_3_15;
    wire logic p_4_16;
    wire logic g_4_16;
    assign p_4_16 = p_3_16 & p_3_8;
    assign g_4_16 = (p_3_16 & g_3_8) | g_3_16;
    wire logic p_4_17;
    wire logic g_4_17;
    assign p_4_17 = p_3_17 & p_3_9;
    assign g_4_17 = (p_3_17 & g_3_9) | g_3_17;
    wire logic p_4_18;
    wire logic g_4_18;
    assign p_4_18 = p_3_18 & p_3_10;
    assign g_4_18 = (p_3_18 & g_3_10) | g_3_18;
    wire logic p_4_19;
    wire logic g_4_19;
    assign p_4_19 = p_3_19 & p_3_11;
    assign g_4_19 = (p_3_19 & g_3_11) | g_3_19;
    wire logic p_4_20;
    wire logic g_4_20;
    assign p_4_20 = p_3_20 & p_3_12;
    assign g_4_20 = (p_3_20 & g_3_12) | g_3_20;
    wire logic p_4_21;
    wire logic g_4_21;
    assign p_4_21 = p_3_21 & p_3_13;
    assign g_4_21 = (p_3_21 & g_3_13) | g_3_21;
    wire logic p_4_22;
    wire logic g_4_22;
    assign p_4_22 = p_3_22 & p_3_14;
    assign g_4_22 = (p_3_22 & g_3_14) | g_3_22;
    wire logic p_4_23;
    wire logic g_4_23;
    assign p_4_23 = p_3_23 & p_3_15;
    assign g_4_23 = (p_3_23 & g_3_15) | g_3_23;
    wire logic p_4_24;
    wire logic g_4_24;
    assign p_4_24 = p_3_24 & p_3_16;
    assign g_4_24 = (p_3_24 & g_3_16) | g_3_24;
    wire logic p_4_25;
    wire logic g_4_25;
    assign p_4_25 = p_3_25 & p_3_17;
    assign g_4_25 = (p_3_25 & g_3_17) | g_3_25;
    wire logic p_4_26;
    wire logic g_4_26;
    assign p_4_26 = p_3_26 & p_3_18;
    assign g_4_26 = (p_3_26 & g_3_18) | g_3_26;
    wire logic p_4_27;
    wire logic g_4_27;
    assign p_4_27 = p_3_27 & p_3_19;
    assign g_4_27 = (p_3_27 & g_3_19) | g_3_27;
    wire logic p_4_28;
    wire logic g_4_28;
    assign p_4_28 = p_3_28 & p_3_20;
    assign g_4_28 = (p_3_28 & g_3_20) | g_3_28;
    wire logic p_4_29;
    wire logic g_4_29;
    assign p_4_29 = p_3_29 & p_3_21;
    assign g_4_29 = (p_3_29 & g_3_21) | g_3_29;
    wire logic p_4_30;
    wire logic g_4_30;
    assign p_4_30 = p_3_30 & p_3_22;
    assign g_4_30 = (p_3_30 & g_3_22) | g_3_30;
    wire logic p_4_31;
    wire logic g_4_31;
    assign p_4_31 = p_3_31 & p_3_23;
    assign g_4_31 = (p_3_31 & g_3_23) | g_3_31;
    
    // KS stage 5
    wire logic p_5_16;
    wire logic g_5_16;
    assign p_5_16 = p_4_16 & p_0[0];
    assign g_5_16 = (p_4_16 & g_0[0]) | g_4_16;
    wire logic p_5_17;
    wire logic g_5_17;
    assign p_5_17 = p_4_17 & p_1_1;
    assign g_5_17 = (p_4_17 & g_1_1) | g_4_17;
    wire logic p_5_18;
    wire logic g_5_18;
    assign p_5_18 = p_4_18 & p_2_2;
    assign g_5_18 = (p_4_18 & g_2_2) | g_4_18;
    wire logic p_5_19;
    wire logic g_5_19;
    assign p_5_19 = p_4_19 & p_2_3;
    assign g_5_19 = (p_4_19 & g_2_3) | g_4_19;
    wire logic p_5_20;
    wire logic g_5_20;
    assign p_5_20 = p_4_20 & p_3_4;
    assign g_5_20 = (p_4_20 & g_3_4) | g_4_20;
    wire logic p_5_21;
    wire logic g_5_21;
    assign p_5_21 = p_4_21 & p_3_5;
    assign g_5_21 = (p_4_21 & g_3_5) | g_4_21;
    wire logic p_5_22;
    wire logic g_5_22;
    assign p_5_22 = p_4_22 & p_3_6;
    assign g_5_22 = (p_4_22 & g_3_6) | g_4_22;
    wire logic p_5_23;
    wire logic g_5_23;
    assign p_5_23 = p_4_23 & p_3_7;
    assign g_5_23 = (p_4_23 & g_3_7) | g_4_23;
    wire logic p_5_24;
    wire logic g_5_24;
    assign p_5_24 = p_4_24 & p_4_8;
    assign g_5_24 = (p_4_24 & g_4_8) | g_4_24;
    wire logic p_5_25;
    wire logic g_5_25;
    assign p_5_25 = p_4_25 & p_4_9;
    assign g_5_25 = (p_4_25 & g_4_9) | g_4_25;
    wire logic p_5_26;
    wire logic g_5_26;
    assign p_5_26 = p_4_26 & p_4_10;
    assign g_5_26 = (p_4_26 & g_4_10) | g_4_26;
    wire logic p_5_27;
    wire logic g_5_27;
    assign p_5_27 = p_4_27 & p_4_11;
    assign g_5_27 = (p_4_27 & g_4_11) | g_4_27;
    wire logic p_5_28;
    wire logic g_5_28;
    assign p_5_28 = p_4_28 & p_4_12;
    assign g_5_28 = (p_4_28 & g_4_12) | g_4_28;
    wire logic p_5_29;
    wire logic g_5_29;
    assign p_5_29 = p_4_29 & p_4_13;
    assign g_5_29 = (p_4_29 & g_4_13) | g_4_29;
    wire logic p_5_30;
    wire logic g_5_30;
    assign p_5_30 = p_4_30 & p_4_14;
    assign g_5_30 = (p_4_30 & g_4_14) | g_4_30;
    wire logic p_5_31;
    wire logic g_5_31;
    assign p_5_31 = p_4_31 & p_4_15;
    assign g_5_31 = (p_4_31 & g_4_15) | g_4_31;
    
    // KS postprocess 
    assign OUT[0] = p_0[0];
    assign OUT[1] = p_0[1] ^ g_0[0];
    assign OUT[2] = p_0[2] ^ g_1_1;
    assign OUT[3] = p_0[3] ^ g_2_2;
    assign OUT[4] = p_0[4] ^ g_2_3;
    assign OUT[5] = p_0[5] ^ g_3_4;
    assign OUT[6] = p_0[6] ^ g_3_5;
    assign OUT[7] = p_0[7] ^ g_3_6;
    assign OUT[8] = p_0[8] ^ g_3_7;
    assign OUT[9] = p_0[9] ^ g_4_8;
    assign OUT[10] = p_0[10] ^ g_4_9;
    assign OUT[11] = p_0[11] ^ g_4_10;
    assign OUT[12] = p_0[12] ^ g_4_11;
    assign OUT[13] = p_0[13] ^ g_4_12;
    assign OUT[14] = p_0[14] ^ g_4_13;
    assign OUT[15] = p_0[15] ^ g_4_14;
    assign OUT[16] = p_0[16] ^ g_4_15;
    assign OUT[17] = p_0[17] ^ g_5_16;
    assign OUT[18] = p_0[18] ^ g_5_17;
    assign OUT[19] = p_0[19] ^ g_5_18;
    assign OUT[20] = p_0[20] ^ g_5_19;
    assign OUT[21] = p_0[21] ^ g_5_20;
    assign OUT[22] = p_0[22] ^ g_5_21;
    assign OUT[23] = p_0[23] ^ g_5_22;
    assign OUT[24] = p_0[24] ^ g_5_23;
    assign OUT[25] = p_0[25] ^ g_5_24;
    assign OUT[26] = p_0[26] ^ g_5_25;
    assign OUT[27] = p_0[27] ^ g_5_26;
    assign OUT[28] = p_0[28] ^ g_5_27;
    assign OUT[29] = p_0[29] ^ g_5_28;
    assign OUT[30] = p_0[30] ^ g_5_29;
    assign OUT[31] = p_0[31] ^ g_5_30;
    assign OUT[32] = g_5_31;
endmodule

module KS_32_spec (
        input logic [31:0] IN1,
        input logic [31:0] IN2,
        output logic adder_correct,
        output logic [32:0] spec_res);
    
    assign spec_res = IN1 + IN2;
    wire [32:0] adder_res;
    KS_32 adder(IN1, IN2, adder_res);
    assign adder_correct = ((spec_res == adder_res) ? 1 : 0);
    
endmodule



module ha (
        input logic a,
        input logic b,
        output logic s,
        output logic c);
    
    assign s = a ^ b;
    assign c = a & b;
endmodule



module fa (
        input logic x,
        input logic y,
        input logic z,
        output logic s,
        output logic c);
    
    assign s = x ^ y ^ z;
    assign c = (x & y) | (x & z) | (y & z);
endmodule


