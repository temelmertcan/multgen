// Note: The license below is based on the template at:
// http://opensource.org/licenses/BSD-3-Clause
// Copyright (C) 2020 Regents of the University of Texas
//All rights reserved.

// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are
// met:

// o Redistributions of source code must retain the above copyright
//   notice, this list of conditions and the following disclaimer.

// o Redistributions in binary form must reproduce the above copyright
//   notice, this list of conditions and the following disclaimer in the
//   documentation and/or other materials provided with the distribution.

// o Neither the name of the copyright holders nor the names of its
//   contributors may be used to endorse or promote products derived
//   from this software without specific prior written permission.

// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
// A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT
// HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
// SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT
// LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
// DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
// THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

// Original Author(s):
// Mertcan Temel         <mert@utexas.edu>

// DO NOT REMOVE:
// This file is generated by Temel's multiplier generator. Download from https://github.com/temelmertcan/multgen.


// Specification module to help understand what the design implements.
module DOT_Product_DT_UB4_LF_4_8x8_plus_10_9to0_spec (
        input logic [3:0][7:0] IN1,
        input logic [3:0][7:0] IN2,
        input logic [9:0] IN3,
        output logic design_is_correct, // is set to 1 iff the output of DOT_Product_DT_UB4_LF_4_8x8_plus_10_9to0  matches its spec
        output logic [9:0] design_res,
        output logic [9:0] spec_res);
    
    assign spec_res = (unsigned'(IN1[0]) * unsigned'(IN2[0])) + 
		      (unsigned'(IN1[1]) * unsigned'(IN2[1])) + 
		      (unsigned'(IN1[2]) * unsigned'(IN2[2])) + 
		      (unsigned'(IN1[3]) * unsigned'(IN2[3])) + 
		      unsigned'(IN3);
    DOT_Product_DT_UB4_LF_4_8x8_plus_10_9to0 dot_product(IN1, IN2, IN3, design_res);
    assign design_is_correct = ((spec_res == design_res) ? 1 : 0);
    
endmodule

module DT_UB4_8x8(
        input logic [7:0] IN1,
        input logic [7:0] IN2,
        output logic [9:0] result0,
        output logic [9:0] result1);
    
    
// Creating Partial Products 

    wire [8:0] mult = {1'b0, IN1};
    wire [8:0] mcand = {1'b0, IN2};
    wire [9:0] mcand_1x;
    wire [9:0] mcand_2x;
    assign mcand_1x = {{1{mcand[8]}},  mcand};
    assign mcand_2x = {{0{mcand[8]}},  mcand, 1'b0};
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[1] mult[0] 1'b0
    wire logic select_0_0, select_e_0, select_2x_0, tcomp0, select_ne_0, select_n2x_0;
    assign select_0_0 =  &{mult[1], mult[0], 1'b0} | ~|{mult[1], mult[0], 1'b0};
    assign select_e_0 = ((~ mult[1]) & (mult[0] ^ 1'b0));
    assign select_ne_0 = mult[1] &  (mult[0] ^ 1'b0);
    assign select_2x_0 = (~ mult[1]) & mult[0] & 1'b0;
    assign select_n2x_0 = mult[1] & (~ mult[0]) & (~ 1'b0);
    reg [9:0] pp_0;
    always @(*) begin
       case (1'b1)
          select_0_0   : pp_0 = 0; 
          select_e_0   : pp_0 = mcand_1x; 
          select_2x_0  : pp_0 = mcand_2x; 
          select_n2x_0 : pp_0 = (~ mcand_2x); 
          select_ne_0  : pp_0 = (~ mcand_1x); 
       endcase 
       pp_0[9] = ~pp_0[9]; // flip the MSB 
    end
    assign tcomp0 =  select_n2x_0 | select_ne_0;
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[3] mult[2] mult[1]
    wire logic select_0_1, select_e_1, select_2x_1, tcomp1, select_ne_1, select_n2x_1;
    assign select_0_1 =  &{mult[3], mult[2], mult[1]} | ~|{mult[3], mult[2], mult[1]};
    assign select_e_1 = ((~ mult[3]) & (mult[2] ^ mult[1]));
    assign select_ne_1 = mult[3] &  (mult[2] ^ mult[1]);
    assign select_2x_1 = (~ mult[3]) & mult[2] & mult[1];
    assign select_n2x_1 = mult[3] & (~ mult[2]) & (~ mult[1]);
    reg [9:0] pp_1;
    always @(*) begin
       case (1'b1)
          select_0_1   : pp_1 = 0; 
          select_e_1   : pp_1 = mcand_1x; 
          select_2x_1  : pp_1 = mcand_2x; 
          select_n2x_1 : pp_1 = (~ mcand_2x); 
          select_ne_1  : pp_1 = (~ mcand_1x); 
       endcase 
       pp_1[9] = ~pp_1[9]; // flip the MSB 
    end
    assign tcomp1 =  select_n2x_1 | select_ne_1;
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[5] mult[4] mult[3]
    wire logic select_0_2, select_e_2, select_2x_2, tcomp2, select_ne_2, select_n2x_2;
    assign select_0_2 =  &{mult[5], mult[4], mult[3]} | ~|{mult[5], mult[4], mult[3]};
    assign select_e_2 = ((~ mult[5]) & (mult[4] ^ mult[3]));
    assign select_ne_2 = mult[5] &  (mult[4] ^ mult[3]);
    assign select_2x_2 = (~ mult[5]) & mult[4] & mult[3];
    assign select_n2x_2 = mult[5] & (~ mult[4]) & (~ mult[3]);
    reg [9:0] pp_2;
    always @(*) begin
       case (1'b1)
          select_0_2   : pp_2 = 0; 
          select_e_2   : pp_2 = mcand_1x; 
          select_2x_2  : pp_2 = mcand_2x; 
          select_n2x_2 : pp_2 = (~ mcand_2x); 
          select_ne_2  : pp_2 = (~ mcand_1x); 
       endcase 
       pp_2[9] = ~pp_2[9]; // flip the MSB 
    end
    assign tcomp2 =  select_n2x_2 | select_ne_2;
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[7] mult[6] mult[5]
    wire logic select_0_3, select_e_3, select_2x_3, tcomp3, select_ne_3, select_n2x_3;
    assign select_0_3 =  &{mult[7], mult[6], mult[5]} | ~|{mult[7], mult[6], mult[5]};
    assign select_e_3 = ((~ mult[7]) & (mult[6] ^ mult[5]));
    assign select_ne_3 = mult[7] &  (mult[6] ^ mult[5]);
    assign select_2x_3 = (~ mult[7]) & mult[6] & mult[5];
    assign select_n2x_3 = mult[7] & (~ mult[6]) & (~ mult[5]);
    reg [9:0] pp_3;
    always @(*) begin
       case (1'b1)
          select_0_3   : pp_3 = 0; 
          select_e_3   : pp_3 = mcand_1x; 
          select_2x_3  : pp_3 = mcand_2x; 
          select_n2x_3 : pp_3 = (~ mcand_2x); 
          select_ne_3  : pp_3 = (~ mcand_1x); 
       endcase 
       pp_3[9] = ~pp_3[9]; // flip the MSB 
    end
    assign tcomp3 =  select_n2x_3 | select_ne_3;
    
    // Booth Radix-4 Partial Products. Multiplier selectors: mult[8] mult[8] mult[7]
    wire logic select_0_4, select_e_4, select_2x_4, tcomp4, select_ne_4, select_n2x_4;
    assign select_0_4 =  &{mult[8], mult[8], mult[7]} | ~|{mult[8], mult[8], mult[7]};
    assign select_e_4 = ((~ mult[8]) & (mult[8] ^ mult[7]));
    assign select_ne_4 = mult[8] &  (mult[8] ^ mult[7]);
    assign select_2x_4 = (~ mult[8]) & mult[8] & mult[7];
    assign select_n2x_4 = mult[8] & (~ mult[8]) & (~ mult[7]);
    reg [9:0] pp_4;
    always @(*) begin
       case (1'b1)
          select_0_4   : pp_4 = 0; 
          select_e_4   : pp_4 = mcand_1x; 
          select_2x_4  : pp_4 = mcand_2x; 
          select_n2x_4 : pp_4 = (~ mcand_2x); 
          select_ne_4  : pp_4 = (~ mcand_1x); 
       endcase 
       pp_4[9] = ~pp_4[9]; // flip the MSB 
    end
    assign tcomp4 =  select_n2x_4 | select_ne_4;
    
    // The values to be summed in the summation tree, from LSB (left) to MSB:
     // pp_0[0] pp_0[1] pp_0[2] pp_0[3] pp_0[4] pp_0[5] pp_0[6] pp_0[7] pp_0[8] pp_0[9]   --      --      --      --      --      --      --      --    
     //   --      --    pp_1[0] pp_1[1] pp_1[2] pp_1[3] pp_1[4] pp_1[5] pp_1[6] pp_1[7] pp_1[8] pp_1[9]   --      --      --      --      --      --    
     //   --      --      --      --    pp_2[0] pp_2[1] pp_2[2] pp_2[3] pp_2[4] pp_2[5] pp_2[6] pp_2[7] pp_2[8] pp_2[9]   --      --      --      --    
     //   --      --      --      --      --      --    pp_3[0] pp_3[1] pp_3[2] pp_3[3] pp_3[4] pp_3[5] pp_3[6] pp_3[7] pp_3[8] pp_3[9]   --      --    
     //   --      --      --      --      --      --      --      --    pp_4[0] pp_4[1] pp_4[2] pp_4[3] pp_4[4] pp_4[5] pp_4[6] pp_4[7] pp_4[8] pp_4[9] 
     // tcomp0    --    tcomp1    --    tcomp2    --    tcomp3    --    tcomp4    --      --      --      --      --      --      --      --      --    
     //   --      --      --      --      --      --      --      --      --      --      --      --      --      --      --      --      --      --    
    
// Creating Summation Tree 

    
    // Dadda Summation Stage 1
    logic s0 ,c0;
    ha ha0 (pp_0[6], pp_1[4], s0, c0);
    logic s1 ,c1;
    ha ha1 (pp_0[7], pp_1[5], s1, c1);
    logic s2 ,c2; 
    fa fa2 (pp_0[8], pp_1[6], pp_2[4], s2, c2);
    logic s3 ,c3;
    ha ha3 (pp_3[2], pp_4[0], s3, c3);
    logic s4 ,c4; 
    fa fa4 (pp_0[9], pp_1[7], pp_2[5], s4, c4);
    logic s5 ,c5;
    ha ha5 (pp_3[3], pp_4[1], s5, c5);
    
    // Dadda Summation Stage 2
    logic s6 ,c6;
    ha ha6 (pp_0[4], pp_1[2], s6, c6);
    logic s7 ,c7;
    ha ha7 (pp_0[5], pp_1[3], s7, c7);
    logic s8 ,c8; 
    fa fa8 (pp_2[2], pp_3[0], tcomp3, s8, c8);
    logic s9 ,c9; 
    fa fa9 (pp_2[3], pp_3[1], c0, s9, c9);
    logic s10 ,c10; 
    fa fa10 (tcomp4, c1, s2, s10, c10);
    logic s11 ,c11; 
    fa fa11 (c2, c3, s4, s11, c11);
    
    // Dadda Summation Stage 3
    logic s12 ,c12;
    ha ha12 (pp_0[2], pp_1[0], s12, c12);
    logic s13 ,c13;
    ha ha13 (pp_0[3], pp_1[1], s13, c13);
    logic s14 ,c14; 
    fa fa14 (pp_2[0], tcomp2, s6, s14, c14);
    logic s15 ,c15; 
    fa fa15 (pp_2[1], c6, s7, s15, c15);
    logic s16 ,c16; 
    fa fa16 (s0, c7, s8, s16, c16);
    logic s17 ,c17; 
    fa fa17 (s1, c8, s9, s17, c17);
    logic s18 ,c18; 
    fa fa18 (s3, c9, s10, s18, c18);
    logic s19 ,c19; 
    fa fa19 (s5, c10, s11, s19, c19);
    
    
    assign result0[9:0] = {c18, c17, c16, c15, c14, c13, c12, tcomp1, pp_0[1], pp_0[0] };
    assign result1[9:0] = {s19, s18, s17, s16, s15, s14, s13, s12, 1'b0, tcomp0 };
endmodule



module DOT_Product_DT_UB4_LF_4_8x8_plus_10_9to0(
        input logic [3:0][7:0] IN1,
        input logic [3:0][7:0] IN2,
        input logic [9:0] IN3,
        output logic [9:0] result);
    
    wire logic [9:0] m0_0;
    wire logic [9:0] m0_1;
    wire logic [9:0] m1_0;
    wire logic [9:0] m1_1;
    wire logic [9:0] m2_0;
    wire logic [9:0] m2_1;
    wire logic [9:0] m3_0;
    wire logic [9:0] m3_1;
    
    DT_UB4_8x8 m0 (IN1[0][7:0], IN2[0][7:0], m0_0, m0_1);
    DT_UB4_8x8 m1 (IN1[1][7:0], IN2[1][7:0], m1_0, m1_1);
    DT_UB4_8x8 m2 (IN1[2][7:0], IN2[2][7:0], m2_0, m2_1);
    DT_UB4_8x8 m3 (IN1[3][7:0], IN2[3][7:0], m3_0, m3_1);
    
    // The values to be summed in the summation tree, from LSB (left) to MSB:
     // m0_0[0] m0_0[1] m0_0[2] m0_0[3] m0_0[4] m0_0[5] m0_0[6] m0_0[7] m0_0[8] m0_0[9] 
     // m0_1[0]   --    m0_1[2] m0_1[3] m0_1[4] m0_1[5] m0_1[6] m0_1[7] m0_1[8] m0_1[9] 
     // m1_0[0] m1_0[1] m1_0[2] m1_0[3] m1_0[4] m1_0[5] m1_0[6] m1_0[7] m1_0[8] m1_0[9] 
     // m1_1[0]   --    m1_1[2] m1_1[3] m1_1[4] m1_1[5] m1_1[6] m1_1[7] m1_1[8] m1_1[9] 
     // m2_0[0] m2_0[1] m2_0[2] m2_0[3] m2_0[4] m2_0[5] m2_0[6] m2_0[7] m2_0[8] m2_0[9] 
     // m2_1[0]   --    m2_1[2] m2_1[3] m2_1[4] m2_1[5] m2_1[6] m2_1[7] m2_1[8] m2_1[9] 
     // m3_0[0] m3_0[1] m3_0[2] m3_0[3] m3_0[4] m3_0[5] m3_0[6] m3_0[7] m3_0[8] m3_0[9] 
     // m3_1[0]   --    m3_1[2] m3_1[3] m3_1[4] m3_1[5] m3_1[6] m3_1[7] m3_1[8] m3_1[9] 
     // IN3[0]  IN3[1]  IN3[2]  IN3[3]  IN3[4]  IN3[5]  IN3[6]  IN3[7]  IN3[8]  IN3[9]  
     //   --      --      --      --      --      --      --      --      --      --    
    
    // Dadda Summation Stage 1
    logic s0 ,c0; 
    fa fa0 (m0_0[0], m0_1[0], m1_0[0], s0, c0);
    logic s1 ,c1;
    ha ha1 (m1_1[0], m2_0[0], s1, c1);
    logic s2 ,c2;
    ha ha2 (m0_0[1], m1_0[1], s2, c2);
    logic s3 ,c3; 
    fa fa3 (m0_0[2], m0_1[2], m1_0[2], s3, c3);
    logic s4 ,c4; 
    fa fa4 (m1_1[2], m2_0[2], m2_1[2], s4, c4);
    logic s5 ,c5; 
    fa fa5 (m0_0[3], m0_1[3], m1_0[3], s5, c5);
    logic s6 ,c6; 
    fa fa6 (m1_1[3], m2_0[3], m2_1[3], s6, c6);
    logic s7 ,c7;
    ha ha7 (m3_0[3], m3_1[3], s7, c7);
    logic s8 ,c8; 
    fa fa8 (m0_0[4], m0_1[4], m1_0[4], s8, c8);
    logic s9 ,c9; 
    fa fa9 (m1_1[4], m2_0[4], m2_1[4], s9, c9);
    logic s10 ,c10; 
    fa fa10 (m3_0[4], m3_1[4], IN3[4], s10, c10);
    logic s11 ,c11; 
    fa fa11 (m0_0[5], m0_1[5], m1_0[5], s11, c11);
    logic s12 ,c12; 
    fa fa12 (m1_1[5], m2_0[5], m2_1[5], s12, c12);
    logic s13 ,c13; 
    fa fa13 (m3_0[5], m3_1[5], IN3[5], s13, c13);
    logic s14 ,c14; 
    fa fa14 (m0_0[6], m0_1[6], m1_0[6], s14, c14);
    logic s15 ,c15; 
    fa fa15 (m1_1[6], m2_0[6], m2_1[6], s15, c15);
    logic s16 ,c16; 
    fa fa16 (m3_0[6], m3_1[6], IN3[6], s16, c16);
    logic s17 ,c17; 
    fa fa17 (m0_0[7], m0_1[7], m1_0[7], s17, c17);
    logic s18 ,c18; 
    fa fa18 (m1_1[7], m2_0[7], m2_1[7], s18, c18);
    logic s19 ,c19; 
    fa fa19 (m3_0[7], m3_1[7], IN3[7], s19, c19);
    logic s20 ,c20; 
    fa fa20 (m0_0[8], m0_1[8], m1_0[8], s20, c20);
    logic s21 ,c21; 
    fa fa21 (m1_1[8], m2_0[8], m2_1[8], s21, c21);
    logic s22 ,c22; 
    fa fa22 (m3_0[8], m3_1[8], IN3[8], s22, c22);
    logic s23 ,c23; 
    fa fa23 (m0_0[9], m0_1[9], m1_0[9], s23, c23);
    logic s24 ,c24; 
    fa fa24 (m1_1[9], m2_0[9], m2_1[9], s24, c24);
    logic s25 ,c25; 
    fa fa25 (m3_0[9], m3_1[9], IN3[9], s25, c25);
    
    // Dadda Summation Stage 2
    logic s26 ,c26; 
    fa fa26 (m2_1[0], m3_0[0], m3_1[0], s26, c26);
    logic s27 ,c27; 
    fa fa27 (m2_0[1], m3_0[1], IN3[1], s27, c27);
    logic s28 ,c28;
    ha ha28 (c0, c1, s28, c28);
    logic s29 ,c29; 
    fa fa29 (m3_0[2], m3_1[2], IN3[2], s29, c29);
    logic s30 ,c30; 
    fa fa30 (c2, s3, s4, s30, c30);
    logic s31 ,c31; 
    fa fa31 (IN3[3], c3, c4, s31, c31);
    logic s32 ,c32; 
    fa fa32 (s5, s6, s7, s32, c32);
    logic s33 ,c33; 
    fa fa33 (c5, c6, c7, s33, c33);
    logic s34 ,c34; 
    fa fa34 (s8, s9, s10, s34, c34);
    logic s35 ,c35; 
    fa fa35 (c8, c9, c10, s35, c35);
    logic s36 ,c36; 
    fa fa36 (s11, s12, s13, s36, c36);
    logic s37 ,c37; 
    fa fa37 (c11, c12, c13, s37, c37);
    logic s38 ,c38; 
    fa fa38 (s14, s15, s16, s38, c38);
    logic s39 ,c39; 
    fa fa39 (c14, c15, c16, s39, c39);
    logic s40 ,c40; 
    fa fa40 (s17, s18, s19, s40, c40);
    logic s41 ,c41; 
    fa fa41 (c17, c18, c19, s41, c41);
    logic s42 ,c42; 
    fa fa42 (s20, s21, s22, s42, c42);
    logic s43 ,c43; 
    fa fa43 (c20, c21, c22, s43, c43);
    logic s44 ,c44; 
    fa fa44 (s23, s24, s25, s44, c44);
    
    // Dadda Summation Stage 3
    logic s45 ,c45;
    ha ha45 (IN3[0], s0, s45, c45);
    logic s46 ,c46; 
    fa fa46 (s2, c26, s27, s46, c46);
    logic s47 ,c47; 
    fa fa47 (c27, c28, s29, s47, c47);
    logic s48 ,c48; 
    fa fa48 (c29, c30, s31, s48, c48);
    logic s49 ,c49; 
    fa fa49 (c31, c32, s33, s49, c49);
    logic s50 ,c50; 
    fa fa50 (c33, c34, s35, s50, c50);
    logic s51 ,c51; 
    fa fa51 (c35, c36, s37, s51, c51);
    logic s52 ,c52; 
    fa fa52 (c37, c38, s39, s52, c52);
    logic s53 ,c53; 
    fa fa53 (c39, c40, s41, s53, c53);
    logic s54 ,c54; 
    fa fa54 (c41, c42, s43, s54, c54);
    
    // Dadda Summation Stage 4
    logic s55 ,c55;
    ha ha55 (s1, s26, s55, c55);
    logic s56 ,c56; 
    fa fa56 (s28, c45, s46, s56, c56);
    logic s57 ,c57; 
    fa fa57 (s30, c46, s47, s57, c57);
    logic s58 ,c58; 
    fa fa58 (s32, c47, s48, s58, c58);
    logic s59 ,c59; 
    fa fa59 (s34, c48, s49, s59, c59);
    logic s60 ,c60; 
    fa fa60 (s36, c49, s50, s60, c60);
    logic s61 ,c61; 
    fa fa61 (s38, c50, s51, s61, c61);
    logic s62 ,c62; 
    fa fa62 (s40, c51, s52, s62, c62);
    logic s63 ,c63; 
    fa fa63 (s42, c52, s53, s63, c63);
    logic s64 ,c64; 
    fa fa64 (s44, c53, s54, s64, c64);
    
    logic [10:0] adder_result;
    LF_10 final_adder ({c63, c62, c61, c60, c59, c58, c57, c56, c55, s45 }, {s64, s63, s62, s61, s60, s59, s58, s57, s56, s55 }, adder_result );
    assign result[9:0] = adder_result[9:0];
    

endmodule

module LF_10 ( 
        input logic [9:0] IN1,
        input logic [9:0] IN2,
        output logic [10:0] OUT);
    
    wire logic [9:0] p_0;
    wire logic [9:0] g_0;
    assign g_0 = IN1 & IN2;
    assign p_0 = IN1 ^ IN2;
    
// Ladner-Fischer Adder 

    
    // LF stage 1
    wire logic p_1_1;
    wire logic g_1_1;
    assign p_1_1 = p_0[1] & p_0[0];
    assign g_1_1 = (p_0[1] & g_0[0]) | g_0[1];
    wire logic p_1_3;
    wire logic g_1_3;
    assign p_1_3 = p_0[3] & p_0[2];
    assign g_1_3 = (p_0[3] & g_0[2]) | g_0[3];
    wire logic p_1_5;
    wire logic g_1_5;
    assign p_1_5 = p_0[5] & p_0[4];
    assign g_1_5 = (p_0[5] & g_0[4]) | g_0[5];
    wire logic p_1_7;
    wire logic g_1_7;
    assign p_1_7 = p_0[7] & p_0[6];
    assign g_1_7 = (p_0[7] & g_0[6]) | g_0[7];
    wire logic p_1_9;
    wire logic g_1_9;
    assign p_1_9 = p_0[9] & p_0[8];
    assign g_1_9 = (p_0[9] & g_0[8]) | g_0[9];
    
    // LF stage 2
    wire logic p_2_2;
    wire logic g_2_2;
    assign p_2_2 = p_0[2] & p_1_1;
    assign g_2_2 = (p_0[2] & g_1_1) | g_0[2];
    wire logic p_2_3;
    wire logic g_2_3;
    assign p_2_3 = p_1_3 & p_1_1;
    assign g_2_3 = (p_1_3 & g_1_1) | g_1_3;
    wire logic p_2_6;
    wire logic g_2_6;
    assign p_2_6 = p_0[6] & p_1_5;
    assign g_2_6 = (p_0[6] & g_1_5) | g_0[6];
    wire logic p_2_7;
    wire logic g_2_7;
    assign p_2_7 = p_1_7 & p_1_5;
    assign g_2_7 = (p_1_7 & g_1_5) | g_1_7;
    
    // LF stage 3
    wire logic p_3_4;
    wire logic g_3_4;
    assign p_3_4 = p_0[4] & p_2_3;
    assign g_3_4 = (p_0[4] & g_2_3) | g_0[4];
    wire logic p_3_5;
    wire logic g_3_5;
    assign p_3_5 = p_1_5 & p_2_3;
    assign g_3_5 = (p_1_5 & g_2_3) | g_1_5;
    wire logic p_3_6;
    wire logic g_3_6;
    assign p_3_6 = p_2_6 & p_2_3;
    assign g_3_6 = (p_2_6 & g_2_3) | g_2_6;
    wire logic p_3_7;
    wire logic g_3_7;
    assign p_3_7 = p_2_7 & p_2_3;
    assign g_3_7 = (p_2_7 & g_2_3) | g_2_7;
    
    // LF stage 4
    wire logic p_4_8;
    wire logic g_4_8;
    assign p_4_8 = p_0[8] & p_3_7;
    assign g_4_8 = (p_0[8] & g_3_7) | g_0[8];
    wire logic p_4_9;
    wire logic g_4_9;
    assign p_4_9 = p_1_9 & p_3_7;
    assign g_4_9 = (p_1_9 & g_3_7) | g_1_9;
    
    // LF postprocess 
    assign OUT[0] = p_0[0];
    assign OUT[1] = p_0[1] ^ g_0[0];
    assign OUT[2] = p_0[2] ^ g_1_1;
    assign OUT[3] = p_0[3] ^ g_2_2;
    assign OUT[4] = p_0[4] ^ g_2_3;
    assign OUT[5] = p_0[5] ^ g_3_4;
    assign OUT[6] = p_0[6] ^ g_3_5;
    assign OUT[7] = p_0[7] ^ g_3_6;
    assign OUT[8] = p_0[8] ^ g_3_7;
    assign OUT[9] = p_0[9] ^ g_4_8;
    assign OUT[10] = g_4_9;
endmodule

module LF_10_spec (
        input logic [9:0] IN1,
        input logic [9:0] IN2,
        output logic adder_correct,
        output logic [10:0] spec_res);
    
    assign spec_res = IN1 + IN2;
    wire [10:0] adder_res;
    LF_10 adder(IN1, IN2, adder_res);
    assign adder_correct = ((spec_res == adder_res) ? 1 : 0);
    
endmodule



module ha (
        input logic a,
        input logic b,
        output logic s,
        output logic c);
    
    assign s = a ^ b;
    assign c = a & b;
endmodule



module fa (
        input logic x,
        input logic y,
        input logic z,
        output logic s,
        output logic c);
    
    assign s = x ^ y ^ z;
    assign c = (x & y) | (x & z) | (y & z);
endmodule


