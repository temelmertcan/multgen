// Note: The license below is based on the template at:
// http://opensource.org/licenses/BSD-3-Clause
// Copyright (C) 2020 Regents of the University of Texas
//All rights reserved.

// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are
// met:

// o Redistributions of source code must retain the above copyright
//   notice, this list of conditions and the following disclaimer.

// o Redistributions in binary form must reproduce the above copyright
//   notice, this list of conditions and the following disclaimer in the
//   documentation and/or other materials provided with the distribution.

// o Neither the name of the copyright holders nor the names of its
//   contributors may be used to endorse or promote products derived
//   from this software without specific prior written permission.

// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR
// A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT
// HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL,
// SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT
// LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE,
// DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
// THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

// Original Author(s):
// Mertcan Temel         <mert@utexas.edu>

// DO NOT REMOVE:
// This file is generated by Temel's multiplier generator. Download from https://github.com/temelmertcan/multgen.


// Specification module to help understand what the design implements.
module Merged_DT_SSP_RP_16x16_spec (
        input logic [15:0] IN1,
        input logic [15:0] IN2,
        output logic design_is_correct, // is set to 1 iff the output of Merged_DT_SSP_RP_16x16  matches its spec.
        output logic [31:0] design_res,
        output logic [31:0] spec_res);
    
    assign spec_res = signed'(IN1) * signed'(IN2);
    Merged_DT_SSP_RP_16x16 mult(IN1, IN2, design_res);
    assign design_is_correct = ((spec_res == design_res) ? 1 : 0);
    
endmodule



module DT_SSP_9x9_32(
        input logic [8:0] IN1,
        input logic [8:0] IN2,
        output logic [31:0] result0,
        output logic [31:0] result1);
    
    
// Creating Partial Products 

    wire logic [8:0] pp0;
    wire logic [8:0] pp1;
    wire logic [8:0] pp2;
    wire logic [8:0] pp3;
    wire logic [8:0] pp4;
    wire logic [8:0] pp5;
    wire logic [8:0] pp6;
    wire logic [8:0] pp7;
    wire logic [8:0] pp8;
    assign pp0 = ({9{IN1[0]}} & IN2) ^ ((1'b1)<<8);
    assign pp1 = ({9{IN1[1]}} & IN2) ^ ((1'b1)<<8);
    assign pp2 = ({9{IN1[2]}} & IN2) ^ ((1'b1)<<8);
    assign pp3 = ({9{IN1[3]}} & IN2) ^ ((1'b1)<<8);
    assign pp4 = ({9{IN1[4]}} & IN2) ^ ((1'b1)<<8);
    assign pp5 = ({9{IN1[5]}} & IN2) ^ ((1'b1)<<8);
    assign pp6 = ({9{IN1[6]}} & IN2) ^ ((1'b1)<<8);
    assign pp7 = ({9{IN1[7]}} & IN2) ^ ((1'b1)<<8);
    assign pp8 = ~({9{IN1[8]}} & IN2) ^ ((1'b1)<<8);
    
    // The values to be summed in the summation tree, from LSB (left) to MSB:
     // pp0[0] pp0[1] pp0[2] pp0[3] pp0[4] pp0[5] pp0[6] pp0[7] pp0[8]   --     --     --     --     --     --     --     --     --   
     //   --   pp1[0] pp1[1] pp1[2] pp1[3] pp1[4] pp1[5] pp1[6] pp1[7] pp1[8]   --     --     --     --     --     --     --     --   
     //   --     --   pp2[0] pp2[1] pp2[2] pp2[3] pp2[4] pp2[5] pp2[6] pp2[7] pp2[8]   --     --     --     --     --     --     --   
     //   --     --     --   pp3[0] pp3[1] pp3[2] pp3[3] pp3[4] pp3[5] pp3[6] pp3[7] pp3[8]   --     --     --     --     --     --   
     //   --     --     --     --   pp4[0] pp4[1] pp4[2] pp4[3] pp4[4] pp4[5] pp4[6] pp4[7] pp4[8]   --     --     --     --     --   
     //   --     --     --     --     --   pp5[0] pp5[1] pp5[2] pp5[3] pp5[4] pp5[5] pp5[6] pp5[7] pp5[8]   --     --     --     --   
     //   --     --     --     --     --     --   pp6[0] pp6[1] pp6[2] pp6[3] pp6[4] pp6[5] pp6[6] pp6[7] pp6[8]   --     --     --   
     //   --     --     --     --     --     --     --   pp7[0] pp7[1] pp7[2] pp7[3] pp7[4] pp7[5] pp7[6] pp7[7] pp7[8]   --     --   
     //   --     --     --     --     --     --     --     --   pp8[0] pp8[1] pp8[2] pp8[3] pp8[4] pp8[5] pp8[6] pp8[7] pp8[8]   --   
     //   --     --     --     --     --     --     --     --     --     --     --     --     --     --     --     --     --     --   
    
// Creating Summation Tree 

    
    // Dadda Summation Stage 1
    logic s0 ,c0;
    ha ha0 (pp0[6], pp1[5], s0, c0);
    logic s1 ,c1; 
    fa fa1 (pp0[7], pp1[6], pp2[5], s1, c1);
    logic s2 ,c2;
    ha ha2 (pp3[4], pp4[3], s2, c2);
    logic s3 ,c3; 
    fa fa3 (pp0[8], pp1[7], pp2[6], s3, c3);
    logic s4 ,c4; 
    fa fa4 (pp3[5], pp4[4], pp5[3], s4, c4);
    logic s5 ,c5;
    ha ha5 (pp6[2], pp7[1], s5, c5);
    logic s6 ,c6; 
    fa fa6 (pp1[8], pp2[7], pp3[6], s6, c6);
    logic s7 ,c7; 
    fa fa7 (pp4[5], pp5[4], pp6[3], s7, c7);
    logic s8 ,c8;
    ha ha8 (pp7[2], pp8[1], s8, c8);
    logic s9 ,c9; 
    fa fa9 (pp2[8], pp3[7], pp4[6], s9, c9);
    logic s10 ,c10; 
    fa fa10 (pp5[5], pp6[4], pp7[3], s10, c10);
    logic s11 ,c11; 
    fa fa11 (pp3[8], pp4[7], pp5[6], s11, c11);
    
    // Dadda Summation Stage 2
    logic s12 ,c12;
    ha ha12 (pp0[4], pp1[3], s12, c12);
    logic s13 ,c13; 
    fa fa13 (pp0[5], pp1[4], pp2[3], s13, c13);
    logic s14 ,c14;
    ha ha14 (pp3[2], pp4[1], s14, c14);
    logic s15 ,c15; 
    fa fa15 (pp2[4], pp3[3], pp4[2], s15, c15);
    logic s16 ,c16; 
    fa fa16 (pp5[1], pp6[0], s0, s16, c16);
    logic s17 ,c17; 
    fa fa17 (pp5[2], pp6[1], pp7[0], s17, c17);
    logic s18 ,c18; 
    fa fa18 (c0, s1, s2, s18, c18);
    logic s19 ,c19; 
    fa fa19 (pp8[0], c1, c2, s19, c19);
    logic s20 ,c20; 
    fa fa20 (s3, s4, s5, s20, c20);
    logic s21 ,c21; 
    fa fa21 (c3, c4, c5, s21, c21);
    logic s22 ,c22; 
    fa fa22 (s6, s7, s8, s22, c22);
    logic s23 ,c23; 
    fa fa23 (pp8[2], c6, c7, s23, c23);
    logic s24 ,c24; 
    fa fa24 (c8, s9, s10, s24, c24);
    logic s25 ,c25; 
    fa fa25 (pp6[5], pp7[4], pp8[3], s25, c25);
    logic s26 ,c26; 
    fa fa26 (c9, c10, s11, s26, c26);
    logic s27 ,c27; 
    fa fa27 (pp4[8], pp5[7], pp6[6], s27, c27);
    logic s28 ,c28; 
    fa fa28 (pp7[5], pp8[4], c11, s28, c28);
    logic s29 ,c29; 
    fa fa29 (pp5[8], pp6[7], pp7[6], s29, c29);
    
    // Dadda Summation Stage 3
    logic s30 ,c30;
    ha ha30 (pp0[3], pp1[2], s30, c30);
    logic s31 ,c31; 
    fa fa31 (pp2[2], pp3[1], pp4[0], s31, c31);
    logic s32 ,c32; 
    fa fa32 (pp5[0], c12, s13, s32, c32);
    logic s33 ,c33; 
    fa fa33 (c13, c14, s15, s33, c33);
    logic s34 ,c34; 
    fa fa34 (c15, c16, s17, s34, c34);
    logic s35 ,c35; 
    fa fa35 (c17, c18, s19, s35, c35);
    logic s36 ,c36; 
    fa fa36 (c19, c20, s21, s36, c36);
    logic s37 ,c37; 
    fa fa37 (c21, c22, s23, s37, c37);
    logic s38 ,c38; 
    fa fa38 (c23, c24, s25, s38, c38);
    logic s39 ,c39; 
    fa fa39 (c25, c26, s27, s39, c39);
    logic s40 ,c40; 
    fa fa40 (pp8[5], c27, c28, s40, c40);
    logic s41 ,c41; 
    fa fa41 (pp6[8], pp7[7], pp8[6], s41, c41);
    
    // Dadda Summation Stage 4
    logic s42 ,c42;
    ha ha42 (pp0[2], pp1[1], s42, c42);
    logic s43 ,c43; 
    fa fa43 (pp2[1], pp3[0], s30, s43, c43);
    logic s44 ,c44; 
    fa fa44 (s12, c30, s31, s44, c44);
    logic s45 ,c45; 
    fa fa45 (s14, c31, s32, s45, c45);
    logic s46 ,c46; 
    fa fa46 (s16, c32, s33, s46, c46);
    logic s47 ,c47; 
    fa fa47 (s18, c33, s34, s47, c47);
    logic s48 ,c48; 
    fa fa48 (s20, c34, s35, s48, c48);
    logic s49 ,c49; 
    fa fa49 (s22, c35, s36, s49, c49);
    logic s50 ,c50; 
    fa fa50 (s24, c36, s37, s50, c50);
    logic s51 ,c51; 
    fa fa51 (s26, c37, s38, s51, c51);
    logic s52 ,c52; 
    fa fa52 (s28, c38, s39, s52, c52);
    logic s53 ,c53; 
    fa fa53 (s29, c39, s40, s53, c53);
    logic s54 ,c54; 
    fa fa54 (c29, c40, s41, s54, c54);
    logic s55 ,c55; 
    fa fa55 (pp7[8], pp8[7], c41, s55, c55);
    
    assign result0[0] = pp0[0];
    assign result1[0] = 1'b0;
    
    assign result0[16:1] = {pp8[8], c54, c53, c52, c51, c50, c49, c48, c47, c46, c45, c44, c43, c42, pp2[0], pp0[1] };
    assign result1[16:1] = {c55, s55, s54, s53, s52, s51, s50, s49, s48, s47, s46, s45, s44, s43, s42, pp1[0] };
    assign result0[17] = 1'b0;
    assign result1[17] = 1'b0;
    assign result0[18] = 1'b0;
    assign result1[18] = 1'b0;
    assign result0[19] = 1'b0;
    assign result1[19] = 1'b0;
    assign result0[20] = 1'b0;
    assign result1[20] = 1'b0;
    assign result0[21] = 1'b0;
    assign result1[21] = 1'b0;
    assign result0[22] = 1'b0;
    assign result1[22] = 1'b0;
    assign result0[23] = 1'b0;
    assign result1[23] = 1'b0;
    assign result0[24] = 1'b0;
    assign result1[24] = 1'b0;
    assign result0[25] = 1'b0;
    assign result1[25] = 1'b0;
    assign result0[26] = 1'b0;
    assign result1[26] = 1'b0;
    assign result0[27] = 1'b0;
    assign result1[27] = 1'b0;
    assign result0[28] = 1'b0;
    assign result1[28] = 1'b0;
    assign result0[29] = 1'b0;
    assign result1[29] = 1'b0;
    assign result0[30] = 1'b0;
    assign result1[30] = 1'b0;
    assign result0[31] = 1'b0;
    assign result1[31] = 1'b0;
endmodule



module Merged_DT_SSP_RP_16x16(
        input logic [15:0] IN1,
        input logic [15:0] IN2,
        output logic [31:0] result);
    wire logic [31:0] m1_0;
    wire logic [31:0] m1_1;
    wire logic [31:0] m2_0;
    wire logic [31:0] m2_1;
    wire logic [31:0] m3_0;
    wire logic [31:0] m3_1;
    wire logic [31:0] m4_0;
    wire logic [31:0] m4_1;
    
    DT_SSP_9x9_32 m1 ({1'b0, IN1[7:0]}, {1'b0, IN2[7:0]}, m1_0, m1_1);
    DT_SSP_9x9_32 m2 ({IN2[15], IN2[15:8]}, {1'b0, IN1[7:0]}, m2_0, m2_1);
    DT_SSP_9x9_32 m3 ({IN1[15], IN1[15:8]}, {1'b0, IN2[7:0]}, m3_0, m3_1);
    DT_SSP_9x9_32 m4 ({IN1[15],IN1[15:8]}, {IN2[15], IN2[15:8]}, m4_0, m4_1);
    
    
    // The values to be summed in the summation tree, from LSB (left) to MSB:
     // m1_0[0]  m1_0[1]  m1_0[2]  m1_0[3]  m1_0[4]  m1_0[5]  m1_0[6]  m1_0[7]  m1_0[8]  m1_0[9]  m1_0[10] m1_0[11] m1_0[12] m1_0[13] m1_0[14] m1_0[15] m1_0[16]   --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     
     //   --     m1_1[1]  m1_1[2]  m1_1[3]  m1_1[4]  m1_1[5]  m1_1[6]  m1_1[7]  m1_1[8]  m1_1[9]  m1_1[10] m1_1[11] m1_1[12] m1_1[13] m1_1[14] m1_1[15] m1_1[16]   --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --     m2_0[0]  m2_0[1]  m2_0[2]  m2_0[3]  m2_0[4]  m2_0[5]  m2_0[6]  m2_0[7]  m2_0[8]  m2_0[9]  m2_0[10] m2_0[11] m2_0[12] m2_0[13] m2_0[14] m2_0[15] m2_0[16]   --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --       --     m2_1[1]  m2_1[2]  m2_1[3]  m2_1[4]  m2_1[5]  m2_1[6]  m2_1[7]  m2_1[8]  m2_1[9]  m2_1[10] m2_1[11] m2_1[12] m2_1[13] m2_1[14] m2_1[15] m2_1[16]   --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --     m3_0[0]  m3_0[1]  m3_0[2]  m3_0[3]  m3_0[4]  m3_0[5]  m3_0[6]  m3_0[7]  m3_0[8]  m3_0[9]  m3_0[10] m3_0[11] m3_0[12] m3_0[13] m3_0[14] m3_0[15] m3_0[16]   --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --       --     m3_1[1]  m3_1[2]  m3_1[3]  m3_1[4]  m3_1[5]  m3_1[6]  m3_1[7]  m3_1[8]  m3_1[9]  m3_1[10] m3_1[11] m3_1[12] m3_1[13] m3_1[14] m3_1[15] m3_1[16]   --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     m4_0[0]  m4_0[1]  m4_0[2]  m4_0[3]  m4_0[4]  m4_0[5]  m4_0[6]  m4_0[7]  m4_0[8]  m4_0[9]  m4_0[10] m4_0[11] m4_0[12] m4_0[13] m4_0[14] m4_0[15] 
     //   --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     m4_1[1]  m4_1[2]  m4_1[3]  m4_1[4]  m4_1[5]  m4_1[6]  m4_1[7]  m4_1[8]  m4_1[9]  m4_1[10] m4_1[11] m4_1[12] m4_1[13] m4_1[14] m4_1[15] 
     //   --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --       --     
     //   --       --       --       --       --       --       --       --       --     1'b1       --       --       --       --       --       --       --     1'b1       --       --       --       --       --       --       --     1'b1     1'b1     1'b1     1'b1     1'b1     1'b1     1'b1     
    
    // Dadda Summation Stage 1
    logic s0 ,c0;
    ha ha0 (m1_0[9], m1_1[9], s0, c0);
    logic s1 ,c1;
    ha ha1 (m1_0[10], m1_1[10], s1, c1);
    logic s2 ,c2;
    ha ha2 (m1_0[11], m1_1[11], s2, c2);
    logic s3 ,c3;
    ha ha3 (m1_0[12], m1_1[12], s3, c3);
    logic s4 ,c4;
    ha ha4 (m1_0[13], m1_1[13], s4, c4);
    logic s5 ,c5;
    ha ha5 (m1_0[14], m1_1[14], s5, c5);
    logic s6 ,c6;
    ha ha6 (m1_0[15], m1_1[15], s6, c6);
    logic s7 ,c7; 
    fa fa7 (m1_0[16], m1_1[16], m2_0[8], s7, c7);
    logic s8 ,c8; 
    fa fa8 (m2_0[9], m2_1[9], m3_0[9], s8, c8);
    logic s9 ,c9;
    ha ha9 (m2_0[10], m2_1[10], s9, c9);
    logic s10 ,c10;
    ha ha10 (m2_0[11], m2_1[11], s10, c10);
    logic s11 ,c11;
    ha ha11 (m2_0[12], m2_1[12], s11, c11);
    logic s12 ,c12;
    ha ha12 (m2_0[13], m2_1[13], s12, c12);
    logic s13 ,c13;
    ha ha13 (m2_0[14], m2_1[14], s13, c13);
    logic s14 ,c14;
    ha ha14 (m2_0[15], m2_1[15], s14, c14);
    logic s15 ,c15;
    ha ha15 (m2_0[16], m2_1[16], s15, c15);
    
    // Dadda Summation Stage 2
    logic s16 ,c16; 
    fa fa16 (m2_0[1], m2_1[1], m3_0[1], s16, c16);
    logic s17 ,c17; 
    fa fa17 (m2_0[2], m2_1[2], m3_0[2], s17, c17);
    logic s18 ,c18;
    ha ha18 (m3_1[2], c0, s18, c18);
    logic s19 ,c19; 
    fa fa19 (m2_0[3], m2_1[3], m3_0[3], s19, c19);
    logic s20 ,c20; 
    fa fa20 (m3_1[3], c1, s2, s20, c20);
    logic s21 ,c21; 
    fa fa21 (m2_0[4], m2_1[4], m3_0[4], s21, c21);
    logic s22 ,c22; 
    fa fa22 (m3_1[4], c2, s3, s22, c22);
    logic s23 ,c23; 
    fa fa23 (m2_0[5], m2_1[5], m3_0[5], s23, c23);
    logic s24 ,c24; 
    fa fa24 (m3_1[5], c3, s4, s24, c24);
    logic s25 ,c25; 
    fa fa25 (m2_0[6], m2_1[6], m3_0[6], s25, c25);
    logic s26 ,c26; 
    fa fa26 (m3_1[6], c4, s5, s26, c26);
    logic s27 ,c27; 
    fa fa27 (m2_0[7], m2_1[7], m3_0[7], s27, c27);
    logic s28 ,c28; 
    fa fa28 (m3_1[7], c5, s6, s28, c28);
    logic s29 ,c29; 
    fa fa29 (m2_1[8], m3_0[8], m3_1[8], s29, c29);
    logic s30 ,c30; 
    fa fa30 (m4_0[0], c6, s7, s30, c30);
    logic s31 ,c31; 
    fa fa31 (m3_1[9], m4_0[1], m4_1[1], s31, c31);
    logic s32 ,c32; 
    fa fa32 (1'b1, c7, s8, s32, c32);
    logic s33 ,c33; 
    fa fa33 (m3_0[10], m3_1[10], m4_0[2], s33, c33);
    logic s34 ,c34; 
    fa fa34 (m4_1[2], c8, s9, s34, c34);
    logic s35 ,c35; 
    fa fa35 (m3_0[11], m3_1[11], m4_0[3], s35, c35);
    logic s36 ,c36; 
    fa fa36 (m4_1[3], c9, s10, s36, c36);
    logic s37 ,c37; 
    fa fa37 (m3_0[12], m3_1[12], m4_0[4], s37, c37);
    logic s38 ,c38; 
    fa fa38 (m4_1[4], c10, s11, s38, c38);
    logic s39 ,c39; 
    fa fa39 (m3_0[13], m3_1[13], m4_0[5], s39, c39);
    logic s40 ,c40; 
    fa fa40 (m4_1[5], c11, s12, s40, c40);
    logic s41 ,c41; 
    fa fa41 (m3_0[14], m3_1[14], m4_0[6], s41, c41);
    logic s42 ,c42; 
    fa fa42 (m4_1[6], c12, s13, s42, c42);
    logic s43 ,c43; 
    fa fa43 (m3_0[15], m3_1[15], m4_0[7], s43, c43);
    logic s44 ,c44; 
    fa fa44 (m4_1[7], c13, s14, s44, c44);
    logic s45 ,c45; 
    fa fa45 (m3_0[16], m3_1[16], m4_0[8], s45, c45);
    logic s46 ,c46; 
    fa fa46 (m4_1[8], c14, s15, s46, c46);
    logic s47 ,c47; 
    fa fa47 (m4_0[9], m4_1[9], 1'b1, s47, c47);
    
    // Dadda Summation Stage 3
    logic s48 ,c48;
    ha ha48 (m1_0[8], m1_1[8], s48, c48);
    logic s49 ,c49; 
    fa fa49 (m3_1[1], 1'b1, s0, s49, c49);
    logic s50 ,c50; 
    fa fa50 (s1, c16, s17, s50, c50);
    logic s51 ,c51; 
    fa fa51 (c17, c18, s19, s51, c51);
    logic s52 ,c52; 
    fa fa52 (c19, c20, s21, s52, c52);
    logic s53 ,c53; 
    fa fa53 (c21, c22, s23, s53, c53);
    logic s54 ,c54; 
    fa fa54 (c23, c24, s25, s54, c54);
    logic s55 ,c55; 
    fa fa55 (c25, c26, s27, s55, c55);
    logic s56 ,c56; 
    fa fa56 (c27, c28, s29, s56, c56);
    logic s57 ,c57; 
    fa fa57 (c29, c30, s31, s57, c57);
    logic s58 ,c58; 
    fa fa58 (c31, c32, s33, s58, c58);
    logic s59 ,c59; 
    fa fa59 (c33, c34, s35, s59, c59);
    logic s60 ,c60; 
    fa fa60 (c35, c36, s37, s60, c60);
    logic s61 ,c61; 
    fa fa61 (c37, c38, s39, s61, c61);
    logic s62 ,c62; 
    fa fa62 (c39, c40, s41, s62, c62);
    logic s63 ,c63; 
    fa fa63 (c41, c42, s43, s63, c63);
    logic s64 ,c64; 
    fa fa64 (c43, c44, s45, s64, c64);
    logic s65 ,c65; 
    fa fa65 (c15, c45, c46, s65, c65);
    logic s66 ,c66; 
    fa fa66 (m4_0[10], m4_1[10], 1'b1, s66, c66);
    logic s67 ,c67;
    ha ha67 (m4_0[11], m4_1[11], s67, c67);
    logic s68 ,c68;
    ha ha68 (m4_0[12], m4_1[12], s68, c68);
    logic s69 ,c69;
    ha ha69 (m4_0[13], m4_1[13], s69, c69);
    logic s70 ,c70;
    ha ha70 (m4_0[14], m4_1[14], s70, c70);
    logic s71 ,c71;
    ha ha71 (m4_0[15], m4_1[15], s71, c71);
    
    // Dadda Summation Stage 4
    logic s72 ,c72;
    ha ha72 (m2_0[0], m3_0[0], s72, c72);
    logic s73 ,c73; 
    fa fa73 (s16, c48, s49, s73, c73);
    logic s74 ,c74; 
    fa fa74 (s18, c49, s50, s74, c74);
    logic s75 ,c75; 
    fa fa75 (s20, c50, s51, s75, c75);
    logic s76 ,c76; 
    fa fa76 (s22, c51, s52, s76, c76);
    logic s77 ,c77; 
    fa fa77 (s24, c52, s53, s77, c77);
    logic s78 ,c78; 
    fa fa78 (s26, c53, s54, s78, c78);
    logic s79 ,c79; 
    fa fa79 (s28, c54, s55, s79, c79);
    logic s80 ,c80; 
    fa fa80 (s30, c55, s56, s80, c80);
    logic s81 ,c81; 
    fa fa81 (s32, c56, s57, s81, c81);
    logic s82 ,c82; 
    fa fa82 (s34, c57, s58, s82, c82);
    logic s83 ,c83; 
    fa fa83 (s36, c58, s59, s83, c83);
    logic s84 ,c84; 
    fa fa84 (s38, c59, s60, s84, c84);
    logic s85 ,c85; 
    fa fa85 (s40, c60, s61, s85, c85);
    logic s86 ,c86; 
    fa fa86 (s42, c61, s62, s86, c86);
    logic s87 ,c87; 
    fa fa87 (s44, c62, s63, s87, c87);
    logic s88 ,c88; 
    fa fa88 (s46, c63, s64, s88, c88);
    logic s89 ,c89; 
    fa fa89 (s47, c64, s65, s89, c89);
    logic s90 ,c90; 
    fa fa90 (c47, c65, s66, s90, c90);
    logic s91 ,c91; 
    fa fa91 (1'b1, c66, s67, s91, c91);
    logic s92 ,c92; 
    fa fa92 (1'b1, c67, s68, s92, c92);
    logic s93 ,c93; 
    fa fa93 (1'b1, c68, s69, s93, c93);
    logic s94 ,c94; 
    fa fa94 (1'b1, c69, s70, s94, c94);
    logic s95 ,c95; 
    fa fa95 (1'b1, c70, s71, s95, c95);
    
    assign result[0] = m1_0[0];
    logic [31:0] adder_result;
    RP_31 final_adder ({c94, c93, c92, c91, c90, c89, c88, c87, c86, c85, c84, c83, c82, c81, c80, c79, c78, c77, c76, c75, c74, c73, c72, s48, m1_0[7], m1_0[6], m1_0[5], m1_0[4], m1_0[3], m1_0[2], m1_0[1] }, {s95, s94, s93, s92, s91, s90, s89, s88, s87, s86, s85, s84, s83, s82, s81, s80, s79, s78, s77, s76, s75, s74, s73, s72, m1_1[7], m1_1[6], m1_1[5], m1_1[4], m1_1[3], m1_1[2], m1_1[1] }, adder_result );
    assign result[31:1] = adder_result[30:0];

endmodule

module RP_31 ( 
        input logic [30:0] IN1,
        input logic [30:0] IN2,
        output logic [31:0] OUT);
    
    logic C0, C1, C2, C3, C4, C5, C6, C7, C8, C9, C10, C11, C12, C13, C14, C15, C16, C17, C18, C19, C20, C21, C22, C23, C24, C25, C26, C27, C28, C29, C30, C31;
    ha m0 (IN1[0], IN2[0], OUT[0], C0);
    fa m1 (IN1[1], IN2[1], C0, OUT[1], C1);
    fa m2 (IN1[2], IN2[2], C1, OUT[2], C2);
    fa m3 (IN1[3], IN2[3], C2, OUT[3], C3);
    fa m4 (IN1[4], IN2[4], C3, OUT[4], C4);
    fa m5 (IN1[5], IN2[5], C4, OUT[5], C5);
    fa m6 (IN1[6], IN2[6], C5, OUT[6], C6);
    fa m7 (IN1[7], IN2[7], C6, OUT[7], C7);
    fa m8 (IN1[8], IN2[8], C7, OUT[8], C8);
    fa m9 (IN1[9], IN2[9], C8, OUT[9], C9);
    fa m10 (IN1[10], IN2[10], C9, OUT[10], C10);
    fa m11 (IN1[11], IN2[11], C10, OUT[11], C11);
    fa m12 (IN1[12], IN2[12], C11, OUT[12], C12);
    fa m13 (IN1[13], IN2[13], C12, OUT[13], C13);
    fa m14 (IN1[14], IN2[14], C13, OUT[14], C14);
    fa m15 (IN1[15], IN2[15], C14, OUT[15], C15);
    fa m16 (IN1[16], IN2[16], C15, OUT[16], C16);
    fa m17 (IN1[17], IN2[17], C16, OUT[17], C17);
    fa m18 (IN1[18], IN2[18], C17, OUT[18], C18);
    fa m19 (IN1[19], IN2[19], C18, OUT[19], C19);
    fa m20 (IN1[20], IN2[20], C19, OUT[20], C20);
    fa m21 (IN1[21], IN2[21], C20, OUT[21], C21);
    fa m22 (IN1[22], IN2[22], C21, OUT[22], C22);
    fa m23 (IN1[23], IN2[23], C22, OUT[23], C23);
    fa m24 (IN1[24], IN2[24], C23, OUT[24], C24);
    fa m25 (IN1[25], IN2[25], C24, OUT[25], C25);
    fa m26 (IN1[26], IN2[26], C25, OUT[26], C26);
    fa m27 (IN1[27], IN2[27], C26, OUT[27], C27);
    fa m28 (IN1[28], IN2[28], C27, OUT[28], C28);
    fa m29 (IN1[29], IN2[29], C28, OUT[29], C29);
    fa m30 (IN1[30], IN2[30], C29, OUT[30], C30);
    assign OUT[31] = C30;

endmodule

module RP_31_spec (
        input logic [30:0] IN1,
        input logic [30:0] IN2,
        output logic adder_correct,
        output logic [31:0] spec_res);
    
    assign spec_res = IN1 + IN2;
    wire [31:0] adder_res;
    RP_31 adder(IN1, IN2, adder_res);
    assign adder_correct = ((spec_res == adder_res) ? 1 : 0);
    
endmodule



module ha (
        input logic a,
        input logic b,
        output logic s,
        output logic c);
    
    assign s = a ^ b;
    assign c = a & b;
endmodule



module fa (
        input logic x,
        input logic y,
        input logic z,
        output logic s,
        output logic c);
    
    assign s = x ^ y ^ z;
    assign c = (x & y) | (x & z) | (y & z);
endmodule


